
// 	Thu May  6 05:24:21 2021
//	vlsi
//	localhost.localdomain

module Softmax (\values[0] , \values[1] , \values[2] , \values[3] , \values[4] , 
    \values[5] , \values[6] , \values[7] , \values[8] , \values[9] , class_out);

output [15:0] class_out;
input [15:0] \values[0] ;
input [15:0] \values[1] ;
input [15:0] \values[2] ;
input [15:0] \values[3] ;
input [15:0] \values[4] ;
input [15:0] \values[5] ;
input [15:0] \values[6] ;
input [15:0] \values[7] ;
input [15:0] \values[8] ;
input [15:0] \values[9] ;
wire spw__n672;
wire spw__n671;
wire spw__n646;
wire spw__n645;
wire spw__n644;
wire spw__n46;
wire spt__n7;
wire spt__n4;
wire spt__n1;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire n_0_0_60;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_0_65;
wire n_0_0_66;
wire n_0_0_67;
wire n_0_0_68;
wire n_0_0_69;
wire n_0_0_70;
wire n_0_0_71;
wire n_0_0_72;
wire n_0_0_73;
wire n_0_0_74;
wire n_0_0_75;
wire n_0_0_76;
wire n_0_0_77;
wire n_0_0_78;
wire n_0_0_79;
wire n_0_0_80;
wire n_0_0_81;
wire n_0_0_82;
wire n_0_0_83;
wire n_0_0_84;
wire n_0_0_85;
wire n_0_0_86;
wire n_0_0_87;
wire n_0_0_88;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_93;
wire n_0_0_94;
wire n_0_0_95;
wire n_0_0_96;
wire n_0_0_97;
wire n_0_0_98;
wire n_0_0_99;
wire n_0_0_100;
wire n_0_0_101;
wire n_0_0_102;
wire n_0_0_103;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_0_110;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_0_113;
wire n_0_0_114;
wire n_0_0_115;
wire n_0_0_116;
wire n_0_0_117;
wire n_0_0_118;
wire n_0_0_119;
wire n_0_0_120;
wire n_0_0_121;
wire n_0_0_122;
wire n_0_0_123;
wire n_0_0_124;
wire n_0_0_125;
wire n_0_0_126;
wire n_0_0_127;
wire n_0_0_128;
wire n_0_0_129;
wire n_0_0_130;
wire n_0_0_131;
wire n_0_0_132;
wire n_0_0_133;
wire n_0_0_134;
wire n_0_0_135;
wire n_0_0_136;
wire n_0_0_137;
wire n_0_0_138;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_144;
wire n_0_0_145;
wire n_0_0_146;
wire n_0_0_147;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_0_153;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_0_188;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_0_207;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_0_224;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_0_248;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_0_253;
wire n_0_0_254;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_0_271;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_0_289;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_0_299;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_0_339;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_0_347;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_0_355;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire n_0_0_360;
wire n_0_0_361;
wire n_0_0_362;
wire n_0_0_363;
wire n_0_0_364;
wire n_0_0_365;
wire n_0_0_366;
wire n_0_0_367;
wire n_0_0_368;
wire n_0_0_369;
wire n_0_0_370;
wire n_0_0_371;
wire n_0_0_372;
wire n_0_0_373;
wire n_0_0_374;
wire n_0_0_375;
wire n_0_0_376;
wire n_0_0_377;
wire n_0_0_378;
wire n_0_0_379;
wire n_0_0_380;
wire n_0_0_381;
wire n_0_0_382;
wire n_0_0_383;
wire n_0_0_384;
wire n_0_0_385;
wire n_0_0_386;
wire n_0_0_387;
wire n_0_0_388;
wire n_0_0_389;
wire n_0_0_390;
wire n_0_0_391;
wire n_0_0_392;
wire n_0_0_393;
wire n_0_0_394;
wire n_0_0_395;
wire n_0_0_396;
wire n_0_0_397;
wire n_0_0_398;
wire n_0_0_399;
wire n_0_0_400;
wire n_0_0_401;
wire n_0_0_402;
wire n_0_0_403;
wire n_0_0_404;
wire n_0_0_405;
wire n_0_0_406;
wire n_0_0_407;
wire n_0_0_408;
wire n_0_0_409;
wire n_0_0_410;
wire n_0_0_411;
wire n_0_0_412;
wire n_0_0_413;
wire n_0_0_414;
wire n_0_0_415;
wire n_0_0_416;
wire n_0_0_417;
wire n_0_0_418;
wire n_0_0_419;
wire n_0_0_420;
wire n_0_0_421;
wire n_0_0_422;
wire n_0_0_423;
wire n_0_0_424;
wire n_0_0_425;
wire n_0_0_426;
wire n_0_0_427;
wire n_0_0_428;
wire n_0_0_429;
wire n_0_0_430;
wire n_0_0_431;
wire n_0_0_432;
wire n_0_0_433;
wire n_0_0_434;
wire n_0_0_435;
wire n_0_0_436;
wire n_0_0_437;
wire n_0_0_438;
wire n_0_0_439;
wire n_0_0_440;
wire n_0_0_441;
wire n_0_0_442;
wire n_0_0_443;
wire n_0_0_444;
wire n_0_0_445;
wire n_0_0_446;
wire n_0_0_447;
wire n_0_0_448;
wire n_0_0_449;
wire n_0_0_450;
wire n_0_0_451;
wire n_0_0_452;
wire n_0_0_453;
wire n_0_0_454;
wire n_0_0_455;
wire n_0_0_456;
wire n_0_0_457;
wire n_0_0_458;
wire n_0_0_459;
wire n_0_0_460;
wire n_0_0_461;
wire n_0_0_462;
wire n_0_0_463;
wire n_0_0_464;
wire n_0_0_465;
wire n_0_0_466;
wire n_0_0_467;
wire n_0_0_468;
wire n_0_0_469;
wire n_0_0_470;
wire n_0_0_471;
wire n_0_0_472;
wire n_0_0_473;
wire n_0_0_474;
wire n_0_0_475;
wire n_0_0_476;
wire n_0_0_477;
wire n_0_0_478;
wire n_0_0_479;
wire n_0_0_480;
wire n_0_0_481;
wire n_0_0_482;
wire n_0_0_483;
wire n_0_0_484;
wire n_0_0_485;
wire n_0_0_486;
wire n_0_0_487;
wire n_0_0_488;
wire n_0_0_489;
wire n_0_0_490;
wire n_0_0_491;
wire n_0_0_492;
wire n_0_0_493;
wire n_0_0_494;
wire n_0_0_495;
wire n_0_0_496;
wire n_0_0_497;
wire n_0_0_498;
wire n_0_0_499;
wire n_0_0_500;
wire n_0_0_501;
wire n_0_0_502;
wire n_0_0_503;
wire n_0_0_504;
wire n_0_0_505;
wire n_0_0_506;
wire n_0_0_507;
wire n_0_0_508;
wire n_0_0_509;
wire n_0_0_510;
wire n_0_0_511;
wire n_0_0_512;
wire n_0_0_513;
wire n_0_0_514;
wire n_0_0_515;
wire n_0_0_516;
wire n_0_0_517;
wire n_0_0_518;
wire n_0_0_519;
wire n_0_0_520;
wire n_0_0_521;
wire n_0_0_522;
wire n_0_0_523;
wire n_0_0_524;
wire n_0_0_525;
wire n_0_0_526;
wire spw__n698;
wire spw__n685;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign class_out[15] = class_out[4];
assign class_out[14] = class_out[4];
assign class_out[13] = class_out[4];
assign class_out[12] = class_out[4];
assign class_out[11] = class_out[4];
assign class_out[10] = class_out[4];
assign class_out[9] = class_out[4];
assign class_out[8] = class_out[4];
assign class_out[7] = class_out[4];
assign class_out[6] = class_out[4];
assign class_out[5] = class_out[4];

INV_X1 i_0_0_531 (.ZN (n_0_0_526), .A (\values[0] [15] ));
INV_X1 i_0_0_530 (.ZN (n_0_0_525), .A (\values[0] [14] ));
INV_X1 i_0_0_529 (.ZN (n_0_0_524), .A (\values[0] [13] ));
INV_X1 i_0_0_528 (.ZN (n_0_0_523), .A (\values[0] [12] ));
INV_X1 i_0_0_527 (.ZN (n_0_0_522), .A (\values[0] [11] ));
INV_X1 i_0_0_526 (.ZN (n_0_0_521), .A (\values[0] [10] ));
INV_X1 i_0_0_525 (.ZN (n_0_0_520), .A (\values[0] [8] ));
INV_X1 i_0_0_524 (.ZN (n_0_0_519), .A (\values[0] [7] ));
INV_X1 i_0_0_523 (.ZN (n_0_0_518), .A (\values[0] [6] ));
INV_X1 i_0_0_522 (.ZN (n_0_0_517), .A (\values[0] [4] ));
INV_X1 i_0_0_521 (.ZN (n_0_0_516), .A (\values[0] [3] ));
INV_X16 i_0_0_520 (.ZN (n_0_0_515), .A (\values[0] [1] ));
INV_X1 i_0_0_519 (.ZN (n_0_0_514), .A (\values[1] [9] ));
INV_X1 i_0_0_518 (.ZN (n_0_0_513), .A (\values[1] [5] ));
INV_X16 i_0_0_517 (.ZN (n_0_0_512), .A (\values[1] [2] ));
INV_X1 i_0_0_516 (.ZN (n_0_0_511), .A (\values[3] [12] ));
INV_X1 i_0_0_515 (.ZN (n_0_0_510), .A (\values[4] [1] ));
INV_X1 i_0_0_514 (.ZN (n_0_0_509), .A (\values[5] [15] ));
INV_X1 i_0_0_513 (.ZN (n_0_0_508), .A (\values[6] [15] ));
INV_X1 i_0_0_512 (.ZN (n_0_0_507), .A (\values[8] [1] ));
INV_X1 i_0_0_511 (.ZN (n_0_0_506), .A (\values[8] [0] ));
NOR2_X1 i_0_0_510 (.ZN (n_0_0_505), .A1 (n_0_0_513), .A2 (\values[0] [5] ));
OAI21_X1 i_0_0_509 (.ZN (n_0_0_504), .A (\values[1] [0] ), .B1 (n_0_0_515), .B2 (\values[1] [1] ));
NAND2_X1 i_0_0_508 (.ZN (n_0_0_503), .A1 (n_0_0_515), .A2 (\values[1] [1] ));
OAI221_X1 i_0_0_507 (.ZN (n_0_0_502), .A (n_0_0_503), .B1 (\values[0] [2] ), .B2 (n_0_0_512)
    , .C1 (n_0_0_504), .C2 (\values[0] [0] ));
NAND2_X1 i_0_0_506 (.ZN (n_0_0_501), .A1 (n_0_0_512), .A2 (\values[0] [2] ));
OAI211_X1 i_0_0_505 (.ZN (n_0_0_500), .A (n_0_0_502), .B (n_0_0_501), .C1 (n_0_0_516), .C2 (\values[1] [3] ));
AOI22_X1 i_0_0_504 (.ZN (n_0_0_499), .A1 (n_0_0_517), .A2 (\values[1] [4] ), .B1 (n_0_0_516), .B2 (\values[1] [3] ));
NOR2_X1 i_0_0_503 (.ZN (n_0_0_498), .A1 (n_0_0_517), .A2 (\values[1] [4] ));
AOI221_X2 i_0_0_502 (.ZN (n_0_0_497), .A (n_0_0_498), .B1 (n_0_0_513), .B2 (\values[0] [5] )
    , .C1 (n_0_0_500), .C2 (n_0_0_499));
OAI22_X1 i_0_0_501 (.ZN (n_0_0_496), .A1 (n_0_0_505), .A2 (n_0_0_497), .B1 (n_0_0_518), .B2 (\values[1] [6] ));
AOI22_X1 i_0_0_500 (.ZN (n_0_0_495), .A1 (n_0_0_519), .A2 (\values[1] [7] ), .B1 (n_0_0_518), .B2 (\values[1] [6] ));
NAND2_X1 i_0_0_499 (.ZN (n_0_0_494), .A1 (n_0_0_496), .A2 (n_0_0_495));
OAI221_X1 i_0_0_498 (.ZN (n_0_0_493), .A (n_0_0_494), .B1 (\values[1] [7] ), .B2 (n_0_0_519)
    , .C1 (n_0_0_520), .C2 (\values[1] [8] ));
NAND2_X1 i_0_0_497 (.ZN (n_0_0_492), .A1 (n_0_0_520), .A2 (\values[1] [8] ));
OAI211_X1 i_0_0_496 (.ZN (n_0_0_491), .A (n_0_0_493), .B (n_0_0_492), .C1 (\values[0] [9] ), .C2 (n_0_0_514));
NAND2_X1 i_0_0_495 (.ZN (n_0_0_490), .A1 (n_0_0_514), .A2 (\values[0] [9] ));
OAI211_X1 i_0_0_494 (.ZN (n_0_0_489), .A (n_0_0_491), .B (n_0_0_490), .C1 (n_0_0_521), .C2 (\values[1] [10] ));
AOI22_X1 i_0_0_493 (.ZN (n_0_0_488), .A1 (n_0_0_522), .A2 (\values[1] [11] ), .B1 (n_0_0_521), .B2 (\values[1] [10] ));
NOR2_X1 i_0_0_492 (.ZN (n_0_0_487), .A1 (n_0_0_523), .A2 (\values[1] [12] ));
AOI21_X1 i_0_0_491 (.ZN (n_0_0_486), .A (n_0_0_487), .B1 (n_0_0_489), .B2 (n_0_0_488));
OAI21_X1 i_0_0_490 (.ZN (n_0_0_485), .A (n_0_0_486), .B1 (\values[1] [11] ), .B2 (n_0_0_522));
AOI22_X1 i_0_0_489 (.ZN (n_0_0_484), .A1 (n_0_0_524), .A2 (\values[1] [13] ), .B1 (n_0_0_523), .B2 (\values[1] [12] ));
OAI22_X1 i_0_0_488 (.ZN (n_0_0_483), .A1 (n_0_0_525), .A2 (\values[1] [14] ), .B1 (n_0_0_524), .B2 (\values[1] [13] ));
AOI21_X1 i_0_0_487 (.ZN (n_0_0_482), .A (n_0_0_483), .B1 (n_0_0_485), .B2 (n_0_0_484));
NOR2_X1 i_0_0_486 (.ZN (n_0_0_481), .A1 (n_0_0_526), .A2 (\values[1] [15] ));
AOI211_X1 i_0_0_485 (.ZN (n_0_0_480), .A (n_0_0_482), .B (n_0_0_481), .C1 (n_0_0_525), .C2 (\values[1] [14] ));
AOI21_X2 i_0_0_484 (.ZN (spw__n46), .A (n_0_0_480), .B1 (\values[1] [15] ), .B2 (n_0_0_526));
INV_X4 i_0_0_483 (.ZN (n_0_0_478), .A (n_0_0_479));
NAND2_X1 i_0_0_482 (.ZN (n_0_0_477), .A1 (n_0_0_521), .A2 (spw__n645));
OAI21_X1 i_0_0_481 (.ZN (n_0_0_476), .A (n_0_0_477), .B1 (spw__n645), .B2 (\values[1] [10] ));
NAND2_X1 i_0_0_480 (.ZN (n_0_0_475), .A1 (\values[2] [10] ), .A2 (n_0_0_476));
NAND2_X1 i_0_0_479 (.ZN (n_0_0_474), .A1 (n_0_0_520), .A2 (spw__n644));
OAI21_X1 i_0_0_478 (.ZN (n_0_0_473), .A (n_0_0_474), .B1 (spw__n644), .B2 (\values[1] [8] ));
NOR2_X1 i_0_0_477 (.ZN (n_0_0_472), .A1 (\values[2] [8] ), .A2 (n_0_0_473));
NAND2_X1 i_0_0_476 (.ZN (n_0_0_471), .A1 (n_0_0_519), .A2 (spw__n644));
OAI21_X1 i_0_0_475 (.ZN (n_0_0_470), .A (n_0_0_471), .B1 (n_0_0_478), .B2 (\values[1] [7] ));
NAND2_X1 i_0_0_474 (.ZN (n_0_0_469), .A1 (n_0_0_518), .A2 (n_0_0_478));
OAI21_X1 i_0_0_473 (.ZN (n_0_0_468), .A (n_0_0_469), .B1 (n_0_0_478), .B2 (\values[1] [6] ));
NAND2_X1 i_0_0_472 (.ZN (n_0_0_467), .A1 (n_0_0_468), .A2 (\values[2] [6] ));
NAND2_X1 i_0_0_471 (.ZN (n_0_0_466), .A1 (n_0_0_515), .A2 (n_0_0_478));
OAI21_X2 i_0_0_470 (.ZN (n_0_0_465), .A (n_0_0_466), .B1 (n_0_0_478), .B2 (\values[1] [1] ));
MUX2_X1 i_0_0_469 (.Z (n_0_0_464), .A (\values[0] [0] ), .B (\values[1] [0] ), .S (n_0_0_479));
INV_X1 i_0_0_468 (.ZN (n_0_0_463), .A (n_0_0_464));
OAI211_X1 i_0_0_467 (.ZN (n_0_0_462), .A (n_0_0_463), .B (\values[2] [0] ), .C1 (\values[2] [1] ), .C2 (n_0_0_465));
NAND2_X1 i_0_0_466 (.ZN (n_0_0_461), .A1 (n_0_0_478), .A2 (\values[0] [2] ));
OAI21_X1 i_0_0_465 (.ZN (n_0_0_460), .A (n_0_0_461), .B1 (n_0_0_478), .B2 (n_0_0_512));
INV_X2 i_0_0_464 (.ZN (n_0_0_459), .A (n_0_0_460));
AOI22_X2 i_0_0_463 (.ZN (n_0_0_458), .A1 (\values[2] [1] ), .A2 (n_0_0_465), .B1 (n_0_0_459), .B2 (\values[2] [2] ));
NAND2_X2 i_0_0_462 (.ZN (n_0_0_457), .A1 (n_0_0_516), .A2 (n_0_0_478));
OAI21_X1 i_0_0_461 (.ZN (n_0_0_456), .A (n_0_0_457), .B1 (n_0_0_478), .B2 (\values[1] [3] ));
OAI22_X1 i_0_0_460 (.ZN (n_0_0_455), .A1 (\values[2] [2] ), .A2 (n_0_0_459), .B1 (n_0_0_456), .B2 (\values[2] [3] ));
AOI21_X1 i_0_0_459 (.ZN (n_0_0_454), .A (n_0_0_455), .B1 (n_0_0_462), .B2 (n_0_0_458));
AOI21_X1 i_0_0_458 (.ZN (n_0_0_453), .A (n_0_0_454), .B1 (n_0_0_456), .B2 (\values[2] [3] ));
NAND2_X1 i_0_0_457 (.ZN (n_0_0_452), .A1 (n_0_0_517), .A2 (n_0_0_478));
OAI21_X1 i_0_0_456 (.ZN (n_0_0_451), .A (n_0_0_452), .B1 (n_0_0_478), .B2 (\values[1] [4] ));
NOR2_X1 i_0_0_455 (.ZN (n_0_0_450), .A1 (\values[2] [4] ), .A2 (n_0_0_451));
NAND2_X1 i_0_0_454 (.ZN (n_0_0_449), .A1 (n_0_0_479), .A2 (n_0_0_513));
OAI21_X1 i_0_0_453 (.ZN (n_0_0_448), .A (n_0_0_449), .B1 (n_0_0_479), .B2 (\values[0] [5] ));
AOI22_X1 i_0_0_452 (.ZN (n_0_0_447), .A1 (\values[2] [4] ), .A2 (n_0_0_451), .B1 (n_0_0_448), .B2 (\values[2] [5] ));
OAI21_X1 i_0_0_451 (.ZN (n_0_0_446), .A (n_0_0_447), .B1 (n_0_0_450), .B2 (n_0_0_453));
OAI221_X1 i_0_0_450 (.ZN (n_0_0_445), .A (n_0_0_446), .B1 (n_0_0_448), .B2 (\values[2] [5] )
    , .C1 (\values[2] [6] ), .C2 (n_0_0_468));
NAND2_X1 i_0_0_449 (.ZN (n_0_0_444), .A1 (n_0_0_467), .A2 (n_0_0_445));
OAI21_X1 i_0_0_448 (.ZN (n_0_0_443), .A (n_0_0_444), .B1 (n_0_0_470), .B2 (\values[2] [7] ));
AOI22_X1 i_0_0_447 (.ZN (n_0_0_442), .A1 (\values[2] [8] ), .A2 (n_0_0_473), .B1 (n_0_0_470), .B2 (\values[2] [7] ));
AOI21_X1 i_0_0_446 (.ZN (n_0_0_441), .A (n_0_0_472), .B1 (n_0_0_443), .B2 (n_0_0_442));
NAND2_X1 i_0_0_445 (.ZN (n_0_0_440), .A1 (spw__n645), .A2 (\values[0] [9] ));
OAI21_X1 i_0_0_444 (.ZN (n_0_0_439), .A (n_0_0_440), .B1 (spw__n645), .B2 (n_0_0_514));
INV_X1 i_0_0_443 (.ZN (n_0_0_438), .A (n_0_0_439));
AOI21_X1 i_0_0_442 (.ZN (n_0_0_437), .A (n_0_0_441), .B1 (n_0_0_438), .B2 (\values[2] [9] ));
OAI22_X1 i_0_0_441 (.ZN (n_0_0_436), .A1 (\values[2] [10] ), .A2 (n_0_0_476), .B1 (n_0_0_438), .B2 (\values[2] [9] ));
OAI21_X1 i_0_0_440 (.ZN (n_0_0_435), .A (n_0_0_475), .B1 (n_0_0_437), .B2 (n_0_0_436));
NAND2_X1 i_0_0_439 (.ZN (n_0_0_434), .A1 (n_0_0_522), .A2 (spw__n645));
OAI21_X1 i_0_0_438 (.ZN (n_0_0_433), .A (n_0_0_434), .B1 (spw__n646), .B2 (\values[1] [11] ));
OAI21_X1 i_0_0_437 (.ZN (n_0_0_432), .A (n_0_0_435), .B1 (n_0_0_433), .B2 (\values[2] [11] ));
NAND2_X1 i_0_0_436 (.ZN (n_0_0_431), .A1 (n_0_0_523), .A2 (spw__n646));
OAI21_X1 i_0_0_435 (.ZN (n_0_0_430), .A (n_0_0_431), .B1 (spw__n646), .B2 (\values[1] [12] ));
AOI22_X1 i_0_0_434 (.ZN (n_0_0_429), .A1 (\values[2] [11] ), .A2 (n_0_0_433), .B1 (n_0_0_430), .B2 (\values[2] [12] ));
NAND2_X1 i_0_0_433 (.ZN (n_0_0_428), .A1 (n_0_0_524), .A2 (spw__n646));
OAI21_X1 i_0_0_432 (.ZN (n_0_0_427), .A (n_0_0_428), .B1 (spw__n646), .B2 (\values[1] [13] ));
OAI22_X1 i_0_0_431 (.ZN (n_0_0_426), .A1 (\values[2] [12] ), .A2 (n_0_0_430), .B1 (n_0_0_427), .B2 (\values[2] [13] ));
AOI21_X1 i_0_0_430 (.ZN (n_0_0_425), .A (n_0_0_426), .B1 (n_0_0_432), .B2 (n_0_0_429));
NAND2_X1 i_0_0_429 (.ZN (n_0_0_424), .A1 (n_0_0_525), .A2 (spw__n646));
OAI21_X1 i_0_0_428 (.ZN (n_0_0_423), .A (n_0_0_424), .B1 (spw__n646), .B2 (\values[1] [14] ));
AOI221_X1 i_0_0_427 (.ZN (n_0_0_422), .A (n_0_0_425), .B1 (n_0_0_423), .B2 (\values[2] [14] )
    , .C1 (\values[2] [13] ), .C2 (n_0_0_427));
NAND2_X1 i_0_0_426 (.ZN (n_0_0_421), .A1 (\values[0] [15] ), .A2 (\values[1] [15] ));
NAND2_X1 i_0_0_425 (.ZN (n_0_0_420), .A1 (n_0_0_421), .A2 (\values[2] [15] ));
OAI21_X1 i_0_0_424 (.ZN (n_0_0_419), .A (n_0_0_420), .B1 (n_0_0_423), .B2 (\values[2] [14] ));
OAI22_X2 i_0_0_423 (.ZN (n_0_0_418), .A1 (n_0_0_419), .A2 (n_0_0_422), .B1 (\values[2] [15] ), .B2 (n_0_0_421));
INV_X4 i_0_0_422 (.ZN (n_0_0_417), .A (n_0_0_418));
NAND2_X1 i_0_0_421 (.ZN (n_0_0_416), .A1 (n_0_0_448), .A2 (n_0_0_417));
OAI21_X1 i_0_0_420 (.ZN (n_0_0_415), .A (n_0_0_416), .B1 (n_0_0_417), .B2 (\values[2] [5] ));
NOR2_X1 i_0_0_419 (.ZN (n_0_0_414), .A1 (n_0_0_415), .A2 (\values[3] [5] ));
NAND2_X1 i_0_0_418 (.ZN (n_0_0_413), .A1 (n_0_0_451), .A2 (n_0_0_417));
OAI21_X1 i_0_0_417 (.ZN (n_0_0_412), .A (n_0_0_413), .B1 (n_0_0_417), .B2 (\values[2] [4] ));
NAND2_X1 i_0_0_416 (.ZN (n_0_0_411), .A1 (n_0_0_456), .A2 (n_0_0_417));
OAI21_X1 i_0_0_415 (.ZN (n_0_0_410), .A (n_0_0_411), .B1 (n_0_0_417), .B2 (\values[2] [3] ));
NAND2_X1 i_0_0_414 (.ZN (n_0_0_409), .A1 (n_0_0_410), .A2 (\values[3] [3] ));
NAND2_X2 i_0_0_413 (.ZN (n_0_0_408), .A1 (n_0_0_465), .A2 (n_0_0_417));
OAI21_X1 i_0_0_412 (.ZN (n_0_0_407), .A (n_0_0_408), .B1 (n_0_0_417), .B2 (\values[2] [1] ));
NAND2_X1 i_0_0_411 (.ZN (n_0_0_406), .A1 (n_0_0_418), .A2 (\values[2] [0] ));
OAI21_X1 i_0_0_410 (.ZN (n_0_0_405), .A (n_0_0_406), .B1 (n_0_0_418), .B2 (n_0_0_463));
OAI21_X1 i_0_0_409 (.ZN (n_0_0_404), .A (\values[3] [0] ), .B1 (n_0_0_407), .B2 (\values[3] [1] ));
NOR2_X1 i_0_0_408 (.ZN (n_0_0_403), .A1 (n_0_0_418), .A2 (n_0_0_459));
AOI21_X1 i_0_0_407 (.ZN (spw__n685), .A (n_0_0_403), .B1 (n_0_0_418), .B2 (\values[2] [2] ));
AOI22_X1 i_0_0_406 (.ZN (n_0_0_401), .A1 (\values[3] [1] ), .A2 (n_0_0_407), .B1 (n_0_0_402), .B2 (\values[3] [2] ));
OAI21_X1 i_0_0_405 (.ZN (n_0_0_400), .A (n_0_0_401), .B1 (n_0_0_404), .B2 (n_0_0_405));
OAI221_X1 i_0_0_404 (.ZN (n_0_0_399), .A (n_0_0_400), .B1 (n_0_0_402), .B2 (\values[3] [2] )
    , .C1 (\values[3] [3] ), .C2 (n_0_0_410));
NAND2_X1 i_0_0_403 (.ZN (n_0_0_398), .A1 (n_0_0_409), .A2 (n_0_0_399));
OAI21_X1 i_0_0_402 (.ZN (n_0_0_397), .A (n_0_0_398), .B1 (n_0_0_412), .B2 (\values[3] [4] ));
AOI22_X1 i_0_0_401 (.ZN (n_0_0_396), .A1 (\values[3] [5] ), .A2 (n_0_0_415), .B1 (n_0_0_412), .B2 (\values[3] [4] ));
AOI21_X1 i_0_0_400 (.ZN (n_0_0_395), .A (n_0_0_414), .B1 (n_0_0_397), .B2 (n_0_0_396));
NAND2_X1 i_0_0_399 (.ZN (n_0_0_394), .A1 (n_0_0_417), .A2 (n_0_0_468));
OAI21_X1 i_0_0_398 (.ZN (n_0_0_393), .A (n_0_0_394), .B1 (n_0_0_417), .B2 (\values[2] [6] ));
AOI21_X1 i_0_0_397 (.ZN (n_0_0_392), .A (n_0_0_395), .B1 (n_0_0_393), .B2 (\values[3] [6] ));
NAND2_X1 i_0_0_396 (.ZN (n_0_0_391), .A1 (n_0_0_417), .A2 (n_0_0_470));
OAI21_X1 i_0_0_395 (.ZN (n_0_0_390), .A (n_0_0_391), .B1 (n_0_0_417), .B2 (\values[2] [7] ));
OAI22_X1 i_0_0_394 (.ZN (n_0_0_389), .A1 (\values[3] [6] ), .A2 (n_0_0_393), .B1 (n_0_0_390), .B2 (\values[3] [7] ));
NAND2_X1 i_0_0_393 (.ZN (n_0_0_388), .A1 (n_0_0_473), .A2 (n_0_0_417));
OAI21_X1 i_0_0_392 (.ZN (n_0_0_387), .A (n_0_0_388), .B1 (n_0_0_417), .B2 (\values[2] [8] ));
AOI22_X1 i_0_0_391 (.ZN (n_0_0_386), .A1 (\values[3] [7] ), .A2 (n_0_0_390), .B1 (n_0_0_387), .B2 (\values[3] [8] ));
OAI21_X2 i_0_0_390 (.ZN (n_0_0_385), .A (n_0_0_386), .B1 (n_0_0_392), .B2 (n_0_0_389));
NAND2_X1 i_0_0_389 (.ZN (n_0_0_384), .A1 (n_0_0_418), .A2 (\values[2] [9] ));
OAI21_X1 i_0_0_388 (.ZN (n_0_0_383), .A (n_0_0_384), .B1 (n_0_0_418), .B2 (n_0_0_438));
INV_X1 i_0_0_387 (.ZN (n_0_0_382), .A (n_0_0_383));
OAI221_X1 i_0_0_386 (.ZN (n_0_0_381), .A (n_0_0_385), .B1 (n_0_0_382), .B2 (\values[3] [9] )
    , .C1 (\values[3] [8] ), .C2 (n_0_0_387));
NAND2_X1 i_0_0_385 (.ZN (n_0_0_380), .A1 (n_0_0_476), .A2 (spw__n671));
OAI21_X1 i_0_0_384 (.ZN (n_0_0_379), .A (n_0_0_380), .B1 (spw__n671), .B2 (\values[2] [10] ));
AOI22_X1 i_0_0_383 (.ZN (n_0_0_378), .A1 (\values[3] [9] ), .A2 (n_0_0_382), .B1 (n_0_0_379), .B2 (\values[3] [10] ));
NAND2_X1 i_0_0_382 (.ZN (n_0_0_377), .A1 (n_0_0_433), .A2 (spw__n671));
OAI21_X1 i_0_0_381 (.ZN (n_0_0_376), .A (n_0_0_377), .B1 (spw__n671), .B2 (\values[2] [11] ));
OAI22_X1 i_0_0_380 (.ZN (n_0_0_375), .A1 (\values[3] [10] ), .A2 (n_0_0_379), .B1 (n_0_0_376), .B2 (\values[3] [11] ));
AOI21_X1 i_0_0_379 (.ZN (n_0_0_374), .A (n_0_0_375), .B1 (n_0_0_381), .B2 (n_0_0_378));
AOI21_X1 i_0_0_378 (.ZN (n_0_0_373), .A (n_0_0_374), .B1 (n_0_0_376), .B2 (\values[3] [11] ));
NAND2_X1 i_0_0_377 (.ZN (n_0_0_372), .A1 (spw__n672), .A2 (n_0_0_430));
NAND2_X1 i_0_0_376 (.ZN (n_0_0_371), .A1 (n_0_0_418), .A2 (\values[2] [12] ));
OAI21_X1 i_0_0_375 (.ZN (n_0_0_370), .A (n_0_0_371), .B1 (n_0_0_418), .B2 (n_0_0_430));
OAI21_X1 i_0_0_374 (.ZN (n_0_0_369), .A (n_0_0_372), .B1 (spw__n672), .B2 (\values[2] [12] ));
NOR2_X1 i_0_0_373 (.ZN (n_0_0_368), .A1 (n_0_0_369), .A2 (\values[3] [12] ));
NAND2_X1 i_0_0_372 (.ZN (n_0_0_367), .A1 (n_0_0_427), .A2 (spw__n672));
OAI21_X1 i_0_0_371 (.ZN (n_0_0_366), .A (n_0_0_367), .B1 (spw__n672), .B2 (\values[2] [13] ));
AOI22_X1 i_0_0_370 (.ZN (n_0_0_365), .A1 (\values[3] [12] ), .A2 (n_0_0_369), .B1 (n_0_0_366), .B2 (\values[3] [13] ));
OAI21_X2 i_0_0_369 (.ZN (n_0_0_364), .A (n_0_0_365), .B1 (n_0_0_368), .B2 (n_0_0_373));
NAND2_X1 i_0_0_368 (.ZN (n_0_0_363), .A1 (n_0_0_423), .A2 (spw__n672));
OAI21_X1 i_0_0_367 (.ZN (n_0_0_362), .A (n_0_0_363), .B1 (spw__n672), .B2 (\values[2] [14] ));
OAI221_X1 i_0_0_366 (.ZN (n_0_0_361), .A (n_0_0_364), .B1 (n_0_0_362), .B2 (\values[3] [14] )
    , .C1 (\values[3] [13] ), .C2 (n_0_0_366));
NAND3_X1 i_0_0_365 (.ZN (n_0_0_360), .A1 (\values[0] [15] ), .A2 (\values[1] [15] ), .A3 (\values[2] [15] ));
INV_X1 i_0_0_364 (.ZN (n_0_0_359), .A (n_0_0_360));
NOR2_X1 i_0_0_363 (.ZN (n_0_0_358), .A1 (n_0_0_360), .A2 (\values[3] [15] ));
AOI21_X1 i_0_0_362 (.ZN (n_0_0_357), .A (n_0_0_358), .B1 (n_0_0_362), .B2 (\values[3] [14] ));
AOI22_X4 i_0_0_361 (.ZN (n_0_0_356), .A1 (n_0_0_361), .A2 (n_0_0_357), .B1 (n_0_0_360), .B2 (\values[3] [15] ));
INV_X4 i_0_0_360 (.ZN (n_0_0_355), .A (n_0_0_356));
NAND2_X1 i_0_0_359 (.ZN (n_0_0_354), .A1 (spw__n698), .A2 (spw__n671));
NOR4_X1 i_0_0_358 (.ZN (n_0_0_353), .A1 (\values[0] [11] ), .A2 (\values[0] [10] )
    , .A3 (\values[0] [9] ), .A4 (\values[0] [8] ));
NOR4_X1 i_0_0_357 (.ZN (n_0_0_352), .A1 (n_0_0_526), .A2 (\values[0] [14] ), .A3 (\values[0] [13] ), .A4 (\values[0] [12] ));
NOR4_X1 i_0_0_356 (.ZN (n_0_0_351), .A1 (\values[0] [3] ), .A2 (\values[0] [2] ), .A3 (\values[0] [1] ), .A4 (\values[0] [0] ));
NOR4_X1 i_0_0_355 (.ZN (n_0_0_350), .A1 (\values[0] [7] ), .A2 (\values[0] [6] ), .A3 (\values[0] [5] ), .A4 (\values[0] [4] ));
AND4_X1 i_0_0_354 (.ZN (n_0_0_349), .A1 (n_0_0_353), .A2 (n_0_0_352), .A3 (n_0_0_351), .A4 (n_0_0_350));
NAND2_X1 i_0_0_353 (.ZN (n_0_0_348), .A1 (spw__n645), .A2 (n_0_0_349));
INV_X1 i_0_0_352 (.ZN (n_0_0_347), .A (n_0_0_348));
NOR2_X1 i_0_0_351 (.ZN (n_0_0_346), .A1 (n_0_0_354), .A2 (n_0_0_348));
INV_X1 i_0_0_350 (.ZN (n_0_0_345), .A (n_0_0_346));
NAND2_X1 i_0_0_349 (.ZN (n_0_0_344), .A1 (\values[3] [15] ), .A2 (n_0_0_359));
NAND2_X1 i_0_0_348 (.ZN (n_0_0_343), .A1 (\values[3] [1] ), .A2 (n_0_0_356));
OAI21_X1 i_0_0_347 (.ZN (n_0_0_342), .A (n_0_0_343), .B1 (n_0_0_356), .B2 (n_0_0_407));
MUX2_X1 i_0_0_346 (.Z (n_0_0_341), .A (n_0_0_405), .B (\values[3] [0] ), .S (n_0_0_356));
AOI21_X1 i_0_0_345 (.ZN (n_0_0_340), .A (n_0_0_341), .B1 (n_0_0_342), .B2 (n_0_0_510));
NAND2_X2 i_0_0_344 (.ZN (n_0_0_339), .A1 (n_0_0_402), .A2 (n_0_0_355));
OAI21_X2 i_0_0_343 (.ZN (n_0_0_338), .A (n_0_0_339), .B1 (n_0_0_355), .B2 (\values[3] [2] ));
AOI22_X1 i_0_0_342 (.ZN (n_0_0_337), .A1 (\values[4] [0] ), .A2 (n_0_0_340), .B1 (n_0_0_338), .B2 (\values[4] [2] ));
OAI21_X1 i_0_0_341 (.ZN (n_0_0_336), .A (n_0_0_337), .B1 (n_0_0_342), .B2 (n_0_0_510));
NAND2_X1 i_0_0_340 (.ZN (n_0_0_335), .A1 (n_0_0_410), .A2 (n_0_0_355));
OAI21_X1 i_0_0_339 (.ZN (n_0_0_334), .A (n_0_0_335), .B1 (n_0_0_355), .B2 (\values[3] [3] ));
OAI221_X1 i_0_0_338 (.ZN (n_0_0_333), .A (n_0_0_336), .B1 (n_0_0_334), .B2 (\values[4] [3] )
    , .C1 (\values[4] [2] ), .C2 (n_0_0_338));
NAND2_X1 i_0_0_337 (.ZN (n_0_0_332), .A1 (n_0_0_412), .A2 (n_0_0_355));
OAI21_X1 i_0_0_336 (.ZN (n_0_0_331), .A (n_0_0_332), .B1 (n_0_0_355), .B2 (\values[3] [4] ));
AOI22_X1 i_0_0_335 (.ZN (n_0_0_330), .A1 (\values[4] [3] ), .A2 (n_0_0_334), .B1 (n_0_0_331), .B2 (\values[4] [4] ));
NAND2_X1 i_0_0_334 (.ZN (n_0_0_329), .A1 (n_0_0_415), .A2 (n_0_0_355));
OAI21_X1 i_0_0_333 (.ZN (n_0_0_328), .A (n_0_0_329), .B1 (n_0_0_355), .B2 (\values[3] [5] ));
OAI22_X1 i_0_0_332 (.ZN (n_0_0_327), .A1 (\values[4] [4] ), .A2 (n_0_0_331), .B1 (n_0_0_328), .B2 (\values[4] [5] ));
AOI21_X1 i_0_0_331 (.ZN (n_0_0_326), .A (n_0_0_327), .B1 (n_0_0_333), .B2 (n_0_0_330));
NAND2_X1 i_0_0_330 (.ZN (n_0_0_325), .A1 (n_0_0_355), .A2 (n_0_0_393));
OAI21_X1 i_0_0_329 (.ZN (n_0_0_324), .A (n_0_0_325), .B1 (n_0_0_355), .B2 (\values[3] [6] ));
AOI221_X1 i_0_0_328 (.ZN (n_0_0_323), .A (n_0_0_326), .B1 (n_0_0_324), .B2 (\values[4] [6] )
    , .C1 (\values[4] [5] ), .C2 (n_0_0_328));
NAND2_X1 i_0_0_327 (.ZN (n_0_0_322), .A1 (n_0_0_390), .A2 (n_0_0_355));
OAI21_X1 i_0_0_326 (.ZN (n_0_0_321), .A (n_0_0_322), .B1 (n_0_0_355), .B2 (\values[3] [7] ));
OAI22_X1 i_0_0_325 (.ZN (n_0_0_320), .A1 (\values[4] [6] ), .A2 (n_0_0_324), .B1 (n_0_0_321), .B2 (\values[4] [7] ));
NOR2_X1 i_0_0_324 (.ZN (n_0_0_319), .A1 (n_0_0_323), .A2 (n_0_0_320));
NAND2_X1 i_0_0_323 (.ZN (n_0_0_318), .A1 (n_0_0_387), .A2 (n_0_0_355));
OAI21_X1 i_0_0_322 (.ZN (n_0_0_317), .A (n_0_0_318), .B1 (n_0_0_355), .B2 (\values[3] [8] ));
AOI221_X2 i_0_0_321 (.ZN (n_0_0_316), .A (n_0_0_319), .B1 (n_0_0_317), .B2 (\values[4] [8] )
    , .C1 (\values[4] [7] ), .C2 (n_0_0_321));
NOR2_X1 i_0_0_320 (.ZN (n_0_0_315), .A1 (n_0_0_356), .A2 (n_0_0_382));
AOI21_X1 i_0_0_319 (.ZN (n_0_0_314), .A (n_0_0_315), .B1 (n_0_0_356), .B2 (\values[3] [9] ));
OAI22_X1 i_0_0_318 (.ZN (n_0_0_313), .A1 (\values[4] [8] ), .A2 (n_0_0_317), .B1 (n_0_0_314), .B2 (\values[4] [9] ));
NAND2_X1 i_0_0_317 (.ZN (n_0_0_312), .A1 (n_0_0_379), .A2 (spw__n698));
OAI21_X1 i_0_0_316 (.ZN (n_0_0_311), .A (n_0_0_312), .B1 (spw__n698), .B2 (\values[3] [10] ));
AOI22_X1 i_0_0_315 (.ZN (n_0_0_310), .A1 (\values[4] [9] ), .A2 (n_0_0_314), .B1 (n_0_0_311), .B2 (\values[4] [10] ));
OAI21_X1 i_0_0_314 (.ZN (n_0_0_309), .A (n_0_0_310), .B1 (n_0_0_316), .B2 (n_0_0_313));
NAND2_X1 i_0_0_313 (.ZN (n_0_0_308), .A1 (n_0_0_376), .A2 (spw__n698));
OAI21_X1 i_0_0_312 (.ZN (n_0_0_307), .A (n_0_0_308), .B1 (spw__n698), .B2 (\values[3] [11] ));
OAI22_X1 i_0_0_311 (.ZN (n_0_0_306), .A1 (\values[4] [10] ), .A2 (n_0_0_311), .B1 (n_0_0_307), .B2 (\values[4] [11] ));
INV_X1 i_0_0_310 (.ZN (n_0_0_305), .A (n_0_0_306));
NAND2_X1 i_0_0_309 (.ZN (n_0_0_304), .A1 (n_0_0_356), .A2 (n_0_0_511));
OAI21_X1 i_0_0_308 (.ZN (n_0_0_303), .A (n_0_0_304), .B1 (n_0_0_356), .B2 (n_0_0_370));
AOI222_X1 i_0_0_307 (.ZN (n_0_0_302), .A1 (n_0_0_309), .A2 (n_0_0_305), .B1 (n_0_0_303)
    , .B2 (\values[4] [12] ), .C1 (\values[4] [11] ), .C2 (n_0_0_307));
NAND2_X1 i_0_0_306 (.ZN (n_0_0_301), .A1 (n_0_0_366), .A2 (spw__n698));
OAI21_X1 i_0_0_305 (.ZN (n_0_0_300), .A (n_0_0_301), .B1 (spw__n698), .B2 (\values[3] [13] ));
OAI22_X1 i_0_0_304 (.ZN (n_0_0_299), .A1 (\values[4] [12] ), .A2 (n_0_0_303), .B1 (n_0_0_300), .B2 (\values[4] [13] ));
NAND2_X1 i_0_0_303 (.ZN (n_0_0_298), .A1 (n_0_0_362), .A2 (spw__n698));
OAI21_X1 i_0_0_302 (.ZN (n_0_0_297), .A (n_0_0_298), .B1 (spw__n698), .B2 (\values[3] [14] ));
AOI22_X1 i_0_0_301 (.ZN (n_0_0_296), .A1 (\values[4] [13] ), .A2 (n_0_0_300), .B1 (n_0_0_297), .B2 (\values[4] [14] ));
OAI21_X1 i_0_0_300 (.ZN (n_0_0_295), .A (n_0_0_296), .B1 (n_0_0_302), .B2 (n_0_0_299));
NAND2_X1 i_0_0_299 (.ZN (n_0_0_294), .A1 (n_0_0_344), .A2 (\values[4] [15] ));
OAI211_X1 i_0_0_298 (.ZN (n_0_0_293), .A (n_0_0_295), .B (n_0_0_294), .C1 (\values[4] [14] ), .C2 (n_0_0_297));
OAI21_X4 i_0_0_297 (.ZN (n_0_0_292), .A (n_0_0_293), .B1 (n_0_0_344), .B2 (\values[4] [15] ));
MUX2_X1 i_0_0_296 (.Z (n_0_0_291), .A (n_0_0_341), .B (\values[4] [0] ), .S (n_0_0_292));
INV_X1 i_0_0_295 (.ZN (n_0_0_290), .A (n_0_0_291));
NAND2_X1 i_0_0_294 (.ZN (n_0_0_289), .A1 (n_0_0_510), .A2 (n_0_0_292));
OAI21_X1 i_0_0_293 (.ZN (n_0_0_288), .A (n_0_0_289), .B1 (n_0_0_292), .B2 (n_0_0_342));
AOI22_X2 i_0_0_292 (.ZN (n_0_0_287), .A1 (\values[5] [0] ), .A2 (n_0_0_290), .B1 (n_0_0_288), .B2 (\values[5] [1] ));
NOR2_X1 i_0_0_291 (.ZN (n_0_0_286), .A1 (n_0_0_338), .A2 (n_0_0_292));
AOI21_X1 i_0_0_290 (.ZN (n_0_0_285), .A (n_0_0_286), .B1 (n_0_0_292), .B2 (\values[4] [2] ));
OAI22_X1 i_0_0_289 (.ZN (n_0_0_284), .A1 (\values[5] [1] ), .A2 (n_0_0_288), .B1 (n_0_0_285), .B2 (\values[5] [2] ));
NOR2_X2 i_0_0_288 (.ZN (n_0_0_283), .A1 (n_0_0_334), .A2 (n_0_0_292));
AOI21_X1 i_0_0_287 (.ZN (n_0_0_282), .A (n_0_0_283), .B1 (n_0_0_292), .B2 (\values[4] [3] ));
AOI22_X1 i_0_0_286 (.ZN (n_0_0_281), .A1 (\values[5] [2] ), .A2 (n_0_0_285), .B1 (n_0_0_282), .B2 (\values[5] [3] ));
OAI21_X1 i_0_0_285 (.ZN (n_0_0_280), .A (n_0_0_281), .B1 (n_0_0_287), .B2 (n_0_0_284));
NOR2_X1 i_0_0_284 (.ZN (n_0_0_279), .A1 (n_0_0_331), .A2 (n_0_0_292));
AOI21_X1 i_0_0_283 (.ZN (n_0_0_278), .A (n_0_0_279), .B1 (n_0_0_292), .B2 (\values[4] [4] ));
OAI221_X1 i_0_0_282 (.ZN (n_0_0_277), .A (n_0_0_280), .B1 (n_0_0_278), .B2 (\values[5] [4] )
    , .C1 (\values[5] [3] ), .C2 (n_0_0_282));
NOR2_X1 i_0_0_281 (.ZN (n_0_0_276), .A1 (n_0_0_328), .A2 (n_0_0_292));
AOI21_X1 i_0_0_280 (.ZN (n_0_0_275), .A (n_0_0_276), .B1 (n_0_0_292), .B2 (\values[4] [5] ));
AOI22_X1 i_0_0_279 (.ZN (n_0_0_274), .A1 (\values[5] [4] ), .A2 (n_0_0_278), .B1 (n_0_0_275), .B2 (\values[5] [5] ));
NOR2_X1 i_0_0_278 (.ZN (n_0_0_273), .A1 (n_0_0_324), .A2 (n_0_0_292));
AOI21_X1 i_0_0_277 (.ZN (n_0_0_272), .A (n_0_0_273), .B1 (n_0_0_292), .B2 (\values[4] [6] ));
OAI22_X1 i_0_0_276 (.ZN (n_0_0_271), .A1 (\values[5] [5] ), .A2 (n_0_0_275), .B1 (n_0_0_272), .B2 (\values[5] [6] ));
AOI21_X2 i_0_0_275 (.ZN (n_0_0_270), .A (n_0_0_271), .B1 (n_0_0_277), .B2 (n_0_0_274));
NOR2_X1 i_0_0_274 (.ZN (n_0_0_269), .A1 (n_0_0_321), .A2 (n_0_0_292));
AOI21_X1 i_0_0_273 (.ZN (n_0_0_268), .A (n_0_0_269), .B1 (n_0_0_292), .B2 (\values[4] [7] ));
AOI221_X2 i_0_0_272 (.ZN (n_0_0_267), .A (n_0_0_270), .B1 (n_0_0_268), .B2 (\values[5] [7] )
    , .C1 (\values[5] [6] ), .C2 (n_0_0_272));
NOR2_X1 i_0_0_271 (.ZN (n_0_0_266), .A1 (n_0_0_317), .A2 (n_0_0_292));
AOI21_X1 i_0_0_270 (.ZN (n_0_0_265), .A (n_0_0_266), .B1 (n_0_0_292), .B2 (\values[4] [8] ));
OAI22_X1 i_0_0_269 (.ZN (n_0_0_264), .A1 (\values[5] [7] ), .A2 (n_0_0_268), .B1 (n_0_0_265), .B2 (\values[5] [8] ));
NOR2_X1 i_0_0_268 (.ZN (n_0_0_263), .A1 (n_0_0_314), .A2 (n_0_0_292));
AOI21_X1 i_0_0_267 (.ZN (n_0_0_262), .A (n_0_0_263), .B1 (n_0_0_292), .B2 (\values[4] [9] ));
AOI22_X1 i_0_0_266 (.ZN (n_0_0_261), .A1 (\values[5] [8] ), .A2 (n_0_0_265), .B1 (n_0_0_262), .B2 (\values[5] [9] ));
OAI21_X1 i_0_0_265 (.ZN (n_0_0_260), .A (n_0_0_261), .B1 (n_0_0_267), .B2 (n_0_0_264));
NOR2_X1 i_0_0_264 (.ZN (n_0_0_259), .A1 (n_0_0_311), .A2 (n_0_0_292));
AOI21_X1 i_0_0_263 (.ZN (n_0_0_258), .A (n_0_0_259), .B1 (n_0_0_292), .B2 (\values[4] [10] ));
OAI221_X1 i_0_0_262 (.ZN (n_0_0_257), .A (n_0_0_260), .B1 (n_0_0_258), .B2 (\values[5] [10] )
    , .C1 (\values[5] [9] ), .C2 (n_0_0_262));
NOR2_X1 i_0_0_261 (.ZN (n_0_0_256), .A1 (n_0_0_307), .A2 (n_0_0_292));
AOI21_X1 i_0_0_260 (.ZN (n_0_0_255), .A (n_0_0_256), .B1 (n_0_0_292), .B2 (\values[4] [11] ));
AOI22_X1 i_0_0_259 (.ZN (n_0_0_254), .A1 (\values[5] [10] ), .A2 (n_0_0_258), .B1 (n_0_0_255), .B2 (\values[5] [11] ));
NOR2_X1 i_0_0_258 (.ZN (n_0_0_253), .A1 (n_0_0_303), .A2 (n_0_0_292));
AOI21_X1 i_0_0_257 (.ZN (n_0_0_252), .A (n_0_0_253), .B1 (n_0_0_292), .B2 (\values[4] [12] ));
OAI22_X1 i_0_0_256 (.ZN (n_0_0_251), .A1 (\values[5] [11] ), .A2 (n_0_0_255), .B1 (n_0_0_252), .B2 (\values[5] [12] ));
AOI21_X1 i_0_0_255 (.ZN (n_0_0_250), .A (n_0_0_251), .B1 (n_0_0_257), .B2 (n_0_0_254));
NOR2_X1 i_0_0_254 (.ZN (n_0_0_249), .A1 (n_0_0_300), .A2 (n_0_0_292));
AOI21_X1 i_0_0_253 (.ZN (n_0_0_248), .A (n_0_0_249), .B1 (n_0_0_292), .B2 (\values[4] [13] ));
AOI221_X1 i_0_0_252 (.ZN (n_0_0_247), .A (n_0_0_250), .B1 (n_0_0_248), .B2 (\values[5] [13] )
    , .C1 (\values[5] [12] ), .C2 (n_0_0_252));
NOR2_X1 i_0_0_251 (.ZN (n_0_0_246), .A1 (n_0_0_297), .A2 (n_0_0_292));
AOI21_X1 i_0_0_250 (.ZN (n_0_0_245), .A (n_0_0_246), .B1 (n_0_0_292), .B2 (\values[4] [14] ));
NOR2_X1 i_0_0_249 (.ZN (n_0_0_244), .A1 (n_0_0_245), .A2 (\values[5] [14] ));
NAND3_X1 i_0_0_248 (.ZN (n_0_0_243), .A1 (\values[3] [15] ), .A2 (\values[4] [15] ), .A3 (n_0_0_359));
INV_X1 i_0_0_247 (.ZN (n_0_0_242), .A (n_0_0_243));
AOI211_X1 i_0_0_246 (.ZN (n_0_0_241), .A (n_0_0_247), .B (n_0_0_244), .C1 (n_0_0_243), .C2 (\values[5] [15] ));
OAI21_X2 i_0_0_245 (.ZN (n_0_0_240), .A (n_0_0_241), .B1 (n_0_0_248), .B2 (\values[5] [13] ));
OAI211_X1 i_0_0_244 (.ZN (n_0_0_239), .A (n_0_0_245), .B (\values[5] [14] ), .C1 (n_0_0_509), .C2 (n_0_0_242));
OAI211_X4 i_0_0_243 (.ZN (n_0_0_238), .A (n_0_0_240), .B (n_0_0_239), .C1 (\values[5] [15] ), .C2 (n_0_0_243));
NOR2_X1 i_0_0_242 (.ZN (n_0_0_237), .A1 (n_0_0_292), .A2 (n_0_0_238));
NOR2_X1 i_0_0_241 (.ZN (n_0_0_236), .A1 (n_0_0_509), .A2 (n_0_0_243));
NOR2_X1 i_0_0_240 (.ZN (n_0_0_235), .A1 (n_0_0_245), .A2 (n_0_0_238));
AOI21_X1 i_0_0_239 (.ZN (n_0_0_234), .A (n_0_0_235), .B1 (n_0_0_238), .B2 (\values[5] [14] ));
NOR2_X1 i_0_0_238 (.ZN (n_0_0_233), .A1 (n_0_0_234), .A2 (\values[6] [14] ));
NAND2_X1 i_0_0_237 (.ZN (n_0_0_232), .A1 (n_0_0_234), .A2 (\values[6] [14] ));
NOR2_X1 i_0_0_236 (.ZN (n_0_0_231), .A1 (n_0_0_248), .A2 (n_0_0_238));
AOI21_X1 i_0_0_235 (.ZN (n_0_0_230), .A (n_0_0_231), .B1 (n_0_0_238), .B2 (\values[5] [13] ));
NOR2_X1 i_0_0_234 (.ZN (n_0_0_229), .A1 (n_0_0_238), .A2 (n_0_0_252));
AOI21_X1 i_0_0_233 (.ZN (n_0_0_228), .A (n_0_0_229), .B1 (n_0_0_238), .B2 (\values[5] [12] ));
NOR2_X1 i_0_0_232 (.ZN (n_0_0_227), .A1 (n_0_0_238), .A2 (n_0_0_285));
AOI21_X1 i_0_0_231 (.ZN (n_0_0_226), .A (n_0_0_227), .B1 (n_0_0_238), .B2 (\values[5] [2] ));
NOR2_X1 i_0_0_230 (.ZN (n_0_0_225), .A1 (n_0_0_238), .A2 (n_0_0_288));
AOI21_X1 i_0_0_229 (.ZN (n_0_0_224), .A (n_0_0_225), .B1 (n_0_0_238), .B2 (\values[5] [1] ));
NAND2_X1 i_0_0_228 (.ZN (n_0_0_223), .A1 (n_0_0_238), .A2 (\values[5] [0] ));
OAI21_X1 i_0_0_227 (.ZN (n_0_0_222), .A (n_0_0_223), .B1 (n_0_0_238), .B2 (n_0_0_290));
INV_X1 i_0_0_226 (.ZN (n_0_0_221), .A (n_0_0_222));
OAI211_X1 i_0_0_225 (.ZN (n_0_0_220), .A (\values[6] [0] ), .B (n_0_0_221), .C1 (n_0_0_224), .C2 (\values[6] [1] ));
AOI22_X2 i_0_0_224 (.ZN (n_0_0_219), .A1 (\values[6] [2] ), .A2 (n_0_0_226), .B1 (n_0_0_224), .B2 (\values[6] [1] ));
NOR2_X1 i_0_0_223 (.ZN (n_0_0_218), .A1 (n_0_0_238), .A2 (n_0_0_282));
AOI21_X1 i_0_0_222 (.ZN (n_0_0_217), .A (n_0_0_218), .B1 (n_0_0_238), .B2 (\values[5] [3] ));
OAI22_X1 i_0_0_221 (.ZN (n_0_0_216), .A1 (\values[6] [2] ), .A2 (n_0_0_226), .B1 (n_0_0_217), .B2 (\values[6] [3] ));
AOI21_X1 i_0_0_220 (.ZN (n_0_0_215), .A (n_0_0_216), .B1 (n_0_0_219), .B2 (n_0_0_220));
NOR2_X1 i_0_0_219 (.ZN (n_0_0_214), .A1 (n_0_0_238), .A2 (n_0_0_278));
AOI21_X1 i_0_0_218 (.ZN (n_0_0_213), .A (n_0_0_214), .B1 (n_0_0_238), .B2 (\values[5] [4] ));
AOI221_X1 i_0_0_217 (.ZN (n_0_0_212), .A (n_0_0_215), .B1 (n_0_0_213), .B2 (\values[6] [4] )
    , .C1 (\values[6] [3] ), .C2 (n_0_0_217));
NOR2_X1 i_0_0_216 (.ZN (n_0_0_211), .A1 (n_0_0_238), .A2 (n_0_0_275));
AOI21_X1 i_0_0_215 (.ZN (n_0_0_210), .A (n_0_0_211), .B1 (n_0_0_238), .B2 (\values[5] [5] ));
OAI22_X1 i_0_0_214 (.ZN (n_0_0_209), .A1 (\values[6] [4] ), .A2 (n_0_0_213), .B1 (n_0_0_210), .B2 (\values[6] [5] ));
NOR2_X1 i_0_0_213 (.ZN (n_0_0_208), .A1 (n_0_0_238), .A2 (n_0_0_272));
AOI21_X1 i_0_0_212 (.ZN (n_0_0_207), .A (n_0_0_208), .B1 (n_0_0_238), .B2 (\values[5] [6] ));
AOI22_X1 i_0_0_211 (.ZN (n_0_0_206), .A1 (\values[6] [5] ), .A2 (n_0_0_210), .B1 (n_0_0_207), .B2 (\values[6] [6] ));
OAI21_X1 i_0_0_210 (.ZN (n_0_0_205), .A (n_0_0_206), .B1 (n_0_0_212), .B2 (n_0_0_209));
NOR2_X1 i_0_0_209 (.ZN (n_0_0_204), .A1 (n_0_0_238), .A2 (n_0_0_268));
AOI21_X1 i_0_0_208 (.ZN (n_0_0_203), .A (n_0_0_204), .B1 (n_0_0_238), .B2 (\values[5] [7] ));
OAI221_X1 i_0_0_207 (.ZN (n_0_0_202), .A (n_0_0_205), .B1 (n_0_0_203), .B2 (\values[6] [7] )
    , .C1 (\values[6] [6] ), .C2 (n_0_0_207));
NOR2_X1 i_0_0_206 (.ZN (n_0_0_201), .A1 (n_0_0_238), .A2 (n_0_0_265));
AOI21_X1 i_0_0_205 (.ZN (n_0_0_200), .A (n_0_0_201), .B1 (n_0_0_238), .B2 (\values[5] [8] ));
AOI22_X1 i_0_0_204 (.ZN (n_0_0_199), .A1 (\values[6] [7] ), .A2 (n_0_0_203), .B1 (n_0_0_200), .B2 (\values[6] [8] ));
NOR2_X1 i_0_0_203 (.ZN (n_0_0_198), .A1 (n_0_0_262), .A2 (n_0_0_238));
AOI21_X1 i_0_0_202 (.ZN (n_0_0_197), .A (n_0_0_198), .B1 (n_0_0_238), .B2 (\values[5] [9] ));
OAI22_X1 i_0_0_201 (.ZN (n_0_0_196), .A1 (\values[6] [8] ), .A2 (n_0_0_200), .B1 (n_0_0_197), .B2 (\values[6] [9] ));
AOI21_X1 i_0_0_200 (.ZN (n_0_0_195), .A (n_0_0_196), .B1 (n_0_0_202), .B2 (n_0_0_199));
NOR2_X1 i_0_0_199 (.ZN (n_0_0_194), .A1 (n_0_0_238), .A2 (n_0_0_258));
AOI21_X1 i_0_0_198 (.ZN (n_0_0_193), .A (n_0_0_194), .B1 (n_0_0_238), .B2 (\values[5] [10] ));
AOI221_X1 i_0_0_197 (.ZN (n_0_0_192), .A (n_0_0_195), .B1 (n_0_0_193), .B2 (\values[6] [10] )
    , .C1 (\values[6] [9] ), .C2 (n_0_0_197));
NOR2_X1 i_0_0_196 (.ZN (n_0_0_191), .A1 (n_0_0_238), .A2 (n_0_0_255));
AOI21_X1 i_0_0_195 (.ZN (n_0_0_190), .A (n_0_0_191), .B1 (n_0_0_238), .B2 (\values[5] [11] ));
NOR2_X1 i_0_0_194 (.ZN (n_0_0_189), .A1 (n_0_0_193), .A2 (\values[6] [10] ));
NAND2_X1 i_0_0_193 (.ZN (n_0_0_188), .A1 (n_0_0_228), .A2 (\values[6] [12] ));
NAND2_X1 i_0_0_192 (.ZN (n_0_0_187), .A1 (n_0_0_190), .A2 (\values[6] [11] ));
OAI21_X1 i_0_0_191 (.ZN (n_0_0_186), .A (n_0_0_187), .B1 (n_0_0_189), .B2 (n_0_0_192));
OAI221_X1 i_0_0_190 (.ZN (n_0_0_185), .A (n_0_0_186), .B1 (n_0_0_190), .B2 (\values[6] [11] )
    , .C1 (\values[6] [12] ), .C2 (n_0_0_228));
NAND2_X1 i_0_0_189 (.ZN (n_0_0_184), .A1 (n_0_0_230), .A2 (\values[6] [13] ));
NAND3_X1 i_0_0_188 (.ZN (n_0_0_183), .A1 (n_0_0_188), .A2 (n_0_0_185), .A3 (n_0_0_184));
OAI21_X1 i_0_0_187 (.ZN (n_0_0_182), .A (n_0_0_183), .B1 (n_0_0_230), .B2 (\values[6] [13] ));
OAI21_X2 i_0_0_186 (.ZN (n_0_0_181), .A (n_0_0_232), .B1 (n_0_0_182), .B2 (n_0_0_233));
AOI21_X1 i_0_0_185 (.ZN (n_0_0_180), .A (n_0_0_508), .B1 (n_0_0_236), .B2 (n_0_0_181));
NOR2_X1 i_0_0_184 (.ZN (n_0_0_179), .A1 (n_0_0_236), .A2 (n_0_0_181));
OR2_X4 i_0_0_183 (.ZN (n_0_0_178), .A1 (n_0_0_180), .A2 (n_0_0_179));
INV_X4 i_0_0_182 (.ZN (n_0_0_177), .A (n_0_0_178));
AND2_X1 i_0_0_181 (.ZN (n_0_0_176), .A1 (\values[6] [15] ), .A2 (n_0_0_236));
NAND2_X1 i_0_0_180 (.ZN (n_0_0_175), .A1 (\values[6] [15] ), .A2 (n_0_0_236));
NAND2_X1 i_0_0_179 (.ZN (n_0_0_174), .A1 (n_0_0_200), .A2 (n_0_0_178));
OAI21_X1 i_0_0_178 (.ZN (n_0_0_173), .A (n_0_0_174), .B1 (n_0_0_178), .B2 (\values[6] [8] ));
NAND2_X1 i_0_0_177 (.ZN (n_0_0_172), .A1 (n_0_0_178), .A2 (n_0_0_217));
OAI21_X1 i_0_0_176 (.ZN (n_0_0_171), .A (n_0_0_172), .B1 (n_0_0_178), .B2 (\values[6] [3] ));
NAND2_X1 i_0_0_175 (.ZN (n_0_0_170), .A1 (n_0_0_226), .A2 (n_0_0_178));
OAI21_X1 i_0_0_174 (.ZN (n_0_0_169), .A (n_0_0_170), .B1 (n_0_0_178), .B2 (\values[6] [2] ));
NAND2_X1 i_0_0_173 (.ZN (n_0_0_168), .A1 (\values[6] [0] ), .A2 (n_0_0_177));
OAI21_X1 i_0_0_172 (.ZN (n_0_0_167), .A (n_0_0_168), .B1 (n_0_0_177), .B2 (n_0_0_221));
INV_X1 i_0_0_171 (.ZN (n_0_0_166), .A (n_0_0_167));
NAND2_X1 i_0_0_170 (.ZN (n_0_0_165), .A1 (n_0_0_178), .A2 (n_0_0_224));
OAI21_X1 i_0_0_169 (.ZN (n_0_0_164), .A (n_0_0_165), .B1 (n_0_0_178), .B2 (\values[6] [1] ));
AOI22_X1 i_0_0_168 (.ZN (n_0_0_163), .A1 (\values[7] [0] ), .A2 (n_0_0_166), .B1 (n_0_0_164), .B2 (\values[7] [1] ));
OAI22_X1 i_0_0_167 (.ZN (n_0_0_162), .A1 (\values[7] [2] ), .A2 (n_0_0_169), .B1 (n_0_0_164), .B2 (\values[7] [1] ));
AOI22_X1 i_0_0_166 (.ZN (n_0_0_161), .A1 (\values[7] [3] ), .A2 (n_0_0_171), .B1 (n_0_0_169), .B2 (\values[7] [2] ));
OAI21_X1 i_0_0_165 (.ZN (n_0_0_160), .A (n_0_0_161), .B1 (n_0_0_163), .B2 (n_0_0_162));
NAND2_X1 i_0_0_164 (.ZN (n_0_0_159), .A1 (n_0_0_178), .A2 (n_0_0_213));
OAI21_X1 i_0_0_163 (.ZN (n_0_0_158), .A (n_0_0_159), .B1 (n_0_0_178), .B2 (\values[6] [4] ));
OAI221_X1 i_0_0_162 (.ZN (n_0_0_157), .A (n_0_0_160), .B1 (n_0_0_158), .B2 (\values[7] [4] )
    , .C1 (\values[7] [3] ), .C2 (n_0_0_171));
NAND2_X1 i_0_0_161 (.ZN (n_0_0_156), .A1 (n_0_0_178), .A2 (n_0_0_210));
OAI21_X1 i_0_0_160 (.ZN (n_0_0_155), .A (n_0_0_156), .B1 (n_0_0_178), .B2 (\values[6] [5] ));
AOI22_X1 i_0_0_159 (.ZN (n_0_0_154), .A1 (\values[7] [4] ), .A2 (n_0_0_158), .B1 (n_0_0_155), .B2 (\values[7] [5] ));
NAND2_X1 i_0_0_158 (.ZN (n_0_0_153), .A1 (n_0_0_157), .A2 (n_0_0_154));
NAND2_X1 i_0_0_157 (.ZN (n_0_0_152), .A1 (n_0_0_178), .A2 (n_0_0_207));
OAI21_X1 i_0_0_156 (.ZN (n_0_0_151), .A (n_0_0_152), .B1 (n_0_0_178), .B2 (\values[6] [6] ));
OAI221_X1 i_0_0_155 (.ZN (n_0_0_150), .A (n_0_0_153), .B1 (n_0_0_151), .B2 (\values[7] [6] )
    , .C1 (\values[7] [5] ), .C2 (n_0_0_155));
NAND2_X1 i_0_0_154 (.ZN (n_0_0_149), .A1 (n_0_0_178), .A2 (n_0_0_203));
OAI21_X1 i_0_0_153 (.ZN (n_0_0_148), .A (n_0_0_149), .B1 (n_0_0_178), .B2 (\values[6] [7] ));
AOI22_X1 i_0_0_152 (.ZN (n_0_0_147), .A1 (\values[7] [6] ), .A2 (n_0_0_151), .B1 (n_0_0_148), .B2 (\values[7] [7] ));
OAI22_X1 i_0_0_151 (.ZN (n_0_0_146), .A1 (\values[7] [8] ), .A2 (n_0_0_173), .B1 (n_0_0_148), .B2 (\values[7] [7] ));
AOI21_X1 i_0_0_150 (.ZN (n_0_0_145), .A (n_0_0_146), .B1 (n_0_0_150), .B2 (n_0_0_147));
AOI21_X1 i_0_0_149 (.ZN (n_0_0_144), .A (n_0_0_145), .B1 (n_0_0_173), .B2 (\values[7] [8] ));
NAND2_X1 i_0_0_148 (.ZN (n_0_0_143), .A1 (n_0_0_197), .A2 (n_0_0_178));
OAI21_X1 i_0_0_147 (.ZN (n_0_0_142), .A (n_0_0_143), .B1 (n_0_0_178), .B2 (\values[6] [9] ));
NOR2_X1 i_0_0_146 (.ZN (n_0_0_141), .A1 (\values[7] [9] ), .A2 (n_0_0_142));
NAND2_X1 i_0_0_145 (.ZN (n_0_0_140), .A1 (n_0_0_193), .A2 (n_0_0_178));
OAI21_X1 i_0_0_144 (.ZN (n_0_0_139), .A (n_0_0_140), .B1 (n_0_0_178), .B2 (\values[6] [10] ));
AOI22_X1 i_0_0_143 (.ZN (n_0_0_138), .A1 (\values[7] [9] ), .A2 (n_0_0_142), .B1 (n_0_0_139), .B2 (\values[7] [10] ));
OAI21_X1 i_0_0_142 (.ZN (n_0_0_137), .A (n_0_0_138), .B1 (n_0_0_141), .B2 (n_0_0_144));
NAND2_X1 i_0_0_141 (.ZN (n_0_0_136), .A1 (n_0_0_190), .A2 (n_0_0_178));
OAI21_X1 i_0_0_140 (.ZN (n_0_0_135), .A (n_0_0_136), .B1 (n_0_0_178), .B2 (\values[6] [11] ));
OAI221_X1 i_0_0_139 (.ZN (n_0_0_134), .A (n_0_0_137), .B1 (n_0_0_135), .B2 (\values[7] [11] )
    , .C1 (\values[7] [10] ), .C2 (n_0_0_139));
NAND2_X1 i_0_0_138 (.ZN (n_0_0_133), .A1 (n_0_0_228), .A2 (n_0_0_178));
OAI21_X1 i_0_0_137 (.ZN (n_0_0_132), .A (n_0_0_133), .B1 (n_0_0_178), .B2 (\values[6] [12] ));
AOI22_X1 i_0_0_136 (.ZN (n_0_0_131), .A1 (\values[7] [11] ), .A2 (n_0_0_135), .B1 (n_0_0_132), .B2 (\values[7] [12] ));
NAND2_X1 i_0_0_135 (.ZN (n_0_0_130), .A1 (n_0_0_230), .A2 (n_0_0_178));
OAI21_X1 i_0_0_134 (.ZN (n_0_0_129), .A (n_0_0_130), .B1 (n_0_0_178), .B2 (\values[6] [13] ));
OAI22_X1 i_0_0_133 (.ZN (n_0_0_128), .A1 (\values[7] [12] ), .A2 (n_0_0_132), .B1 (n_0_0_129), .B2 (\values[7] [13] ));
AOI21_X2 i_0_0_132 (.ZN (n_0_0_127), .A (n_0_0_128), .B1 (n_0_0_134), .B2 (n_0_0_131));
NAND2_X1 i_0_0_131 (.ZN (n_0_0_126), .A1 (n_0_0_234), .A2 (n_0_0_178));
OAI21_X1 i_0_0_130 (.ZN (n_0_0_125), .A (n_0_0_126), .B1 (n_0_0_178), .B2 (\values[6] [14] ));
AOI221_X1 i_0_0_129 (.ZN (n_0_0_124), .A (n_0_0_127), .B1 (n_0_0_125), .B2 (\values[7] [14] )
    , .C1 (\values[7] [13] ), .C2 (n_0_0_129));
NAND2_X1 i_0_0_128 (.ZN (n_0_0_123), .A1 (n_0_0_175), .A2 (\values[7] [15] ));
OAI21_X1 i_0_0_127 (.ZN (n_0_0_122), .A (n_0_0_123), .B1 (n_0_0_125), .B2 (\values[7] [14] ));
OAI22_X2 i_0_0_126 (.ZN (spt__n7), .A1 (n_0_0_122), .A2 (n_0_0_124), .B1 (n_0_0_175), .B2 (\values[7] [15] ));
NOR2_X1 i_0_0_125 (.ZN (n_0_0_120), .A1 (n_0_0_121), .A2 (n_0_0_177));
AND2_X1 i_0_0_124 (.ZN (n_0_0_119), .A1 (n_0_0_237), .A2 (n_0_0_120));
NAND2_X1 i_0_0_123 (.ZN (n_0_0_118), .A1 (n_0_0_346), .A2 (n_0_0_119));
NAND2_X2 i_0_0_122 (.ZN (n_0_0_117), .A1 (n_0_0_121), .A2 (\values[7] [1] ));
OAI21_X2 i_0_0_121 (.ZN (n_0_0_116), .A (n_0_0_117), .B1 (n_0_0_121), .B2 (n_0_0_164));
NAND2_X2 i_0_0_120 (.ZN (n_0_0_115), .A1 (n_0_0_121), .A2 (\values[7] [0] ));
OAI21_X1 i_0_0_119 (.ZN (n_0_0_114), .A (n_0_0_115), .B1 (n_0_0_121), .B2 (n_0_0_166));
OAI22_X1 i_0_0_118 (.ZN (n_0_0_113), .A1 (n_0_0_507), .A2 (n_0_0_116), .B1 (n_0_0_114), .B2 (n_0_0_506));
NOR2_X1 i_0_0_117 (.ZN (n_0_0_112), .A1 (n_0_0_121), .A2 (n_0_0_169));
AOI21_X1 i_0_0_116 (.ZN (n_0_0_111), .A (n_0_0_112), .B1 (n_0_0_121), .B2 (\values[7] [2] ));
NAND2_X1 i_0_0_115 (.ZN (n_0_0_110), .A1 (n_0_0_116), .A2 (n_0_0_507));
OAI211_X1 i_0_0_114 (.ZN (n_0_0_109), .A (n_0_0_113), .B (n_0_0_110), .C1 (n_0_0_111), .C2 (\values[8] [2] ));
NOR2_X1 i_0_0_113 (.ZN (n_0_0_108), .A1 (n_0_0_121), .A2 (n_0_0_171));
AOI21_X1 i_0_0_112 (.ZN (n_0_0_107), .A (n_0_0_108), .B1 (n_0_0_121), .B2 (\values[7] [3] ));
AOI22_X2 i_0_0_111 (.ZN (n_0_0_106), .A1 (\values[8] [2] ), .A2 (n_0_0_111), .B1 (n_0_0_107), .B2 (\values[8] [3] ));
NOR2_X1 i_0_0_110 (.ZN (n_0_0_105), .A1 (n_0_0_121), .A2 (n_0_0_158));
AOI21_X1 i_0_0_109 (.ZN (n_0_0_104), .A (n_0_0_105), .B1 (n_0_0_121), .B2 (\values[7] [4] ));
OAI22_X1 i_0_0_108 (.ZN (n_0_0_103), .A1 (\values[8] [3] ), .A2 (n_0_0_107), .B1 (n_0_0_104), .B2 (\values[8] [4] ));
AOI21_X2 i_0_0_107 (.ZN (n_0_0_102), .A (n_0_0_103), .B1 (n_0_0_109), .B2 (n_0_0_106));
NOR2_X1 i_0_0_106 (.ZN (n_0_0_101), .A1 (n_0_0_121), .A2 (n_0_0_155));
AOI21_X1 i_0_0_105 (.ZN (n_0_0_100), .A (n_0_0_101), .B1 (n_0_0_121), .B2 (\values[7] [5] ));
AOI221_X2 i_0_0_104 (.ZN (n_0_0_99), .A (n_0_0_102), .B1 (n_0_0_100), .B2 (\values[8] [5] )
    , .C1 (\values[8] [4] ), .C2 (n_0_0_104));
NOR2_X1 i_0_0_103 (.ZN (n_0_0_98), .A1 (n_0_0_121), .A2 (n_0_0_151));
AOI21_X1 i_0_0_102 (.ZN (n_0_0_97), .A (n_0_0_98), .B1 (n_0_0_121), .B2 (\values[7] [6] ));
OAI22_X1 i_0_0_101 (.ZN (n_0_0_96), .A1 (\values[8] [5] ), .A2 (n_0_0_100), .B1 (n_0_0_97), .B2 (\values[8] [6] ));
NOR2_X1 i_0_0_100 (.ZN (n_0_0_95), .A1 (n_0_0_121), .A2 (n_0_0_148));
AOI21_X1 i_0_0_99 (.ZN (n_0_0_94), .A (n_0_0_95), .B1 (n_0_0_121), .B2 (\values[7] [7] ));
AOI22_X1 i_0_0_98 (.ZN (n_0_0_93), .A1 (\values[8] [6] ), .A2 (n_0_0_97), .B1 (n_0_0_94), .B2 (\values[8] [7] ));
OAI21_X1 i_0_0_97 (.ZN (n_0_0_92), .A (n_0_0_93), .B1 (n_0_0_99), .B2 (n_0_0_96));
NOR2_X1 i_0_0_96 (.ZN (n_0_0_91), .A1 (n_0_0_121), .A2 (n_0_0_173));
AOI21_X1 i_0_0_95 (.ZN (n_0_0_90), .A (n_0_0_91), .B1 (n_0_0_121), .B2 (\values[7] [8] ));
OAI221_X1 i_0_0_94 (.ZN (n_0_0_89), .A (n_0_0_92), .B1 (n_0_0_90), .B2 (\values[8] [8] )
    , .C1 (\values[8] [7] ), .C2 (n_0_0_94));
NOR2_X1 i_0_0_93 (.ZN (n_0_0_88), .A1 (n_0_0_121), .A2 (n_0_0_142));
AOI21_X1 i_0_0_92 (.ZN (n_0_0_87), .A (n_0_0_88), .B1 (n_0_0_121), .B2 (\values[7] [9] ));
AOI22_X1 i_0_0_91 (.ZN (n_0_0_86), .A1 (\values[8] [8] ), .A2 (n_0_0_90), .B1 (n_0_0_87), .B2 (\values[8] [9] ));
NOR2_X1 i_0_0_90 (.ZN (n_0_0_85), .A1 (n_0_0_121), .A2 (n_0_0_139));
AOI21_X1 i_0_0_89 (.ZN (n_0_0_84), .A (n_0_0_85), .B1 (n_0_0_121), .B2 (\values[7] [10] ));
OAI22_X1 i_0_0_88 (.ZN (n_0_0_83), .A1 (\values[8] [9] ), .A2 (n_0_0_87), .B1 (n_0_0_84), .B2 (\values[8] [10] ));
AOI21_X2 i_0_0_87 (.ZN (n_0_0_82), .A (n_0_0_83), .B1 (n_0_0_89), .B2 (n_0_0_86));
NOR2_X1 i_0_0_86 (.ZN (n_0_0_81), .A1 (n_0_0_121), .A2 (n_0_0_135));
AOI21_X1 i_0_0_85 (.ZN (n_0_0_80), .A (n_0_0_81), .B1 (n_0_0_121), .B2 (\values[7] [11] ));
AOI221_X2 i_0_0_84 (.ZN (n_0_0_79), .A (n_0_0_82), .B1 (n_0_0_80), .B2 (\values[8] [11] )
    , .C1 (\values[8] [10] ), .C2 (n_0_0_84));
NOR2_X1 i_0_0_83 (.ZN (n_0_0_78), .A1 (n_0_0_121), .A2 (n_0_0_132));
AOI21_X1 i_0_0_82 (.ZN (n_0_0_77), .A (n_0_0_78), .B1 (n_0_0_121), .B2 (\values[7] [12] ));
OAI22_X1 i_0_0_81 (.ZN (n_0_0_76), .A1 (\values[8] [11] ), .A2 (n_0_0_80), .B1 (n_0_0_77), .B2 (\values[8] [12] ));
NOR2_X1 i_0_0_80 (.ZN (n_0_0_75), .A1 (n_0_0_121), .A2 (n_0_0_129));
AOI21_X1 i_0_0_79 (.ZN (n_0_0_74), .A (n_0_0_75), .B1 (n_0_0_121), .B2 (\values[7] [13] ));
AOI22_X1 i_0_0_78 (.ZN (n_0_0_73), .A1 (\values[8] [12] ), .A2 (n_0_0_77), .B1 (n_0_0_74), .B2 (\values[8] [13] ));
OAI21_X1 i_0_0_77 (.ZN (n_0_0_72), .A (n_0_0_73), .B1 (n_0_0_79), .B2 (n_0_0_76));
NOR2_X1 i_0_0_76 (.ZN (n_0_0_71), .A1 (n_0_0_121), .A2 (n_0_0_125));
AOI21_X1 i_0_0_75 (.ZN (n_0_0_70), .A (n_0_0_71), .B1 (n_0_0_121), .B2 (\values[7] [14] ));
OAI221_X1 i_0_0_74 (.ZN (n_0_0_69), .A (n_0_0_72), .B1 (n_0_0_70), .B2 (\values[8] [14] )
    , .C1 (\values[8] [13] ), .C2 (n_0_0_74));
NAND2_X1 i_0_0_73 (.ZN (n_0_0_68), .A1 (\values[7] [15] ), .A2 (n_0_0_176));
NAND2_X1 i_0_0_72 (.ZN (n_0_0_67), .A1 (n_0_0_70), .A2 (\values[8] [14] ));
OAI211_X2 i_0_0_71 (.ZN (n_0_0_66), .A (n_0_0_69), .B (n_0_0_67), .C1 (n_0_0_68), .C2 (\values[8] [15] ));
NAND2_X1 i_0_0_70 (.ZN (n_0_0_65), .A1 (n_0_0_68), .A2 (\values[8] [15] ));
NAND2_X2 i_0_0_69 (.ZN (spt__n1), .A1 (n_0_0_66), .A2 (n_0_0_65));
NAND3_X1 i_0_0_68 (.ZN (n_0_0_63), .A1 (\values[7] [15] ), .A2 (\values[8] [15] ), .A3 (n_0_0_176));
NAND2_X1 i_0_0_67 (.ZN (n_0_0_62), .A1 (n_0_0_64), .A2 (n_0_0_116));
OAI21_X1 i_0_0_66 (.ZN (n_0_0_61), .A (n_0_0_62), .B1 (n_0_0_64), .B2 (n_0_0_507));
INV_X2 i_0_0_65 (.ZN (n_0_0_60), .A (n_0_0_61));
AND2_X1 i_0_0_64 (.ZN (n_0_0_59), .A1 (n_0_0_114), .A2 (n_0_0_64));
OAI221_X1 i_0_0_63 (.ZN (n_0_0_58), .A (\values[9] [0] ), .B1 (n_0_0_64), .B2 (n_0_0_506)
    , .C1 (n_0_0_60), .C2 (\values[9] [1] ));
NAND2_X1 i_0_0_62 (.ZN (n_0_0_57), .A1 (n_0_0_111), .A2 (n_0_0_64));
OAI21_X1 i_0_0_61 (.ZN (n_0_0_56), .A (n_0_0_57), .B1 (n_0_0_64), .B2 (\values[8] [2] ));
AOI22_X2 i_0_0_60 (.ZN (n_0_0_55), .A1 (\values[9] [1] ), .A2 (n_0_0_60), .B1 (n_0_0_56), .B2 (\values[9] [2] ));
OAI21_X1 i_0_0_59 (.ZN (n_0_0_54), .A (n_0_0_55), .B1 (n_0_0_58), .B2 (n_0_0_59));
NAND2_X1 i_0_0_58 (.ZN (n_0_0_53), .A1 (n_0_0_107), .A2 (n_0_0_64));
OAI21_X1 i_0_0_57 (.ZN (n_0_0_52), .A (n_0_0_53), .B1 (n_0_0_64), .B2 (\values[8] [3] ));
OAI221_X1 i_0_0_56 (.ZN (n_0_0_51), .A (n_0_0_54), .B1 (n_0_0_52), .B2 (\values[9] [3] )
    , .C1 (\values[9] [2] ), .C2 (n_0_0_56));
NAND2_X1 i_0_0_55 (.ZN (n_0_0_50), .A1 (n_0_0_104), .A2 (n_0_0_64));
OAI21_X1 i_0_0_54 (.ZN (n_0_0_49), .A (n_0_0_50), .B1 (n_0_0_64), .B2 (\values[8] [4] ));
AOI22_X1 i_0_0_53 (.ZN (n_0_0_48), .A1 (\values[9] [3] ), .A2 (n_0_0_52), .B1 (n_0_0_49), .B2 (\values[9] [4] ));
NAND2_X1 i_0_0_52 (.ZN (n_0_0_47), .A1 (n_0_0_100), .A2 (n_0_0_64));
OAI21_X1 i_0_0_51 (.ZN (n_0_0_46), .A (n_0_0_47), .B1 (n_0_0_64), .B2 (\values[8] [5] ));
OAI22_X1 i_0_0_50 (.ZN (n_0_0_45), .A1 (\values[9] [4] ), .A2 (n_0_0_49), .B1 (n_0_0_46), .B2 (\values[9] [5] ));
AOI21_X2 i_0_0_49 (.ZN (n_0_0_44), .A (n_0_0_45), .B1 (n_0_0_51), .B2 (n_0_0_48));
NOR2_X1 i_0_0_48 (.ZN (n_0_0_43), .A1 (n_0_0_64), .A2 (\values[8] [6] ));
AOI21_X1 i_0_0_47 (.ZN (n_0_0_42), .A (n_0_0_43), .B1 (n_0_0_64), .B2 (n_0_0_97));
INV_X1 i_0_0_46 (.ZN (n_0_0_41), .A (n_0_0_42));
AOI221_X2 i_0_0_45 (.ZN (n_0_0_40), .A (n_0_0_44), .B1 (n_0_0_41), .B2 (\values[9] [6] )
    , .C1 (\values[9] [5] ), .C2 (n_0_0_46));
NAND2_X1 i_0_0_44 (.ZN (n_0_0_39), .A1 (n_0_0_94), .A2 (n_0_0_64));
OAI21_X1 i_0_0_43 (.ZN (n_0_0_38), .A (n_0_0_39), .B1 (n_0_0_64), .B2 (\values[8] [7] ));
OAI22_X1 i_0_0_42 (.ZN (n_0_0_37), .A1 (\values[9] [6] ), .A2 (n_0_0_41), .B1 (n_0_0_38), .B2 (\values[9] [7] ));
NAND2_X1 i_0_0_41 (.ZN (n_0_0_36), .A1 (n_0_0_90), .A2 (n_0_0_64));
OAI21_X1 i_0_0_40 (.ZN (n_0_0_35), .A (n_0_0_36), .B1 (n_0_0_64), .B2 (\values[8] [8] ));
AOI22_X1 i_0_0_39 (.ZN (n_0_0_34), .A1 (\values[9] [7] ), .A2 (n_0_0_38), .B1 (n_0_0_35), .B2 (\values[9] [8] ));
OAI21_X1 i_0_0_38 (.ZN (n_0_0_33), .A (n_0_0_34), .B1 (n_0_0_40), .B2 (n_0_0_37));
NAND2_X1 i_0_0_37 (.ZN (n_0_0_32), .A1 (n_0_0_87), .A2 (n_0_0_64));
OAI21_X1 i_0_0_36 (.ZN (n_0_0_31), .A (n_0_0_32), .B1 (n_0_0_64), .B2 (\values[8] [9] ));
OAI221_X1 i_0_0_35 (.ZN (n_0_0_30), .A (n_0_0_33), .B1 (n_0_0_31), .B2 (\values[9] [9] )
    , .C1 (\values[9] [8] ), .C2 (n_0_0_35));
NAND2_X1 i_0_0_34 (.ZN (n_0_0_29), .A1 (n_0_0_84), .A2 (n_0_0_64));
OAI21_X1 i_0_0_33 (.ZN (n_0_0_28), .A (n_0_0_29), .B1 (n_0_0_64), .B2 (\values[8] [10] ));
AOI22_X1 i_0_0_32 (.ZN (n_0_0_27), .A1 (\values[9] [9] ), .A2 (n_0_0_31), .B1 (n_0_0_28), .B2 (\values[9] [10] ));
NAND2_X1 i_0_0_31 (.ZN (n_0_0_26), .A1 (n_0_0_80), .A2 (n_0_0_64));
OAI21_X1 i_0_0_30 (.ZN (n_0_0_25), .A (n_0_0_26), .B1 (n_0_0_64), .B2 (\values[8] [11] ));
OAI22_X1 i_0_0_29 (.ZN (n_0_0_24), .A1 (\values[9] [10] ), .A2 (n_0_0_28), .B1 (n_0_0_25), .B2 (\values[9] [11] ));
AOI21_X2 i_0_0_28 (.ZN (n_0_0_23), .A (n_0_0_24), .B1 (n_0_0_30), .B2 (n_0_0_27));
NAND2_X1 i_0_0_27 (.ZN (n_0_0_22), .A1 (n_0_0_77), .A2 (n_0_0_64));
OAI21_X1 i_0_0_26 (.ZN (n_0_0_21), .A (n_0_0_22), .B1 (n_0_0_64), .B2 (\values[8] [12] ));
AOI221_X2 i_0_0_25 (.ZN (n_0_0_20), .A (n_0_0_23), .B1 (n_0_0_21), .B2 (\values[9] [12] )
    , .C1 (\values[9] [11] ), .C2 (n_0_0_25));
NAND2_X1 i_0_0_24 (.ZN (n_0_0_19), .A1 (n_0_0_74), .A2 (n_0_0_64));
OAI21_X1 i_0_0_23 (.ZN (n_0_0_18), .A (n_0_0_19), .B1 (n_0_0_64), .B2 (\values[8] [13] ));
OAI22_X1 i_0_0_22 (.ZN (n_0_0_17), .A1 (\values[9] [12] ), .A2 (n_0_0_21), .B1 (n_0_0_18), .B2 (\values[9] [13] ));
NAND2_X1 i_0_0_21 (.ZN (n_0_0_16), .A1 (\values[9] [13] ), .A2 (n_0_0_18));
OAI21_X1 i_0_0_20 (.ZN (n_0_0_15), .A (n_0_0_16), .B1 (n_0_0_20), .B2 (n_0_0_17));
NAND2_X1 i_0_0_19 (.ZN (n_0_0_14), .A1 (n_0_0_70), .A2 (n_0_0_64));
OAI21_X1 i_0_0_18 (.ZN (n_0_0_13), .A (n_0_0_14), .B1 (n_0_0_64), .B2 (\values[8] [14] ));
OAI21_X1 i_0_0_17 (.ZN (n_0_0_12), .A (n_0_0_15), .B1 (n_0_0_13), .B2 (\values[9] [14] ));
NOR2_X1 i_0_0_16 (.ZN (n_0_0_11), .A1 (n_0_0_63), .A2 (\values[9] [15] ));
AOI21_X1 i_0_0_15 (.ZN (n_0_0_10), .A (n_0_0_11), .B1 (n_0_0_13), .B2 (\values[9] [14] ));
AOI22_X1 i_0_0_14 (.ZN (n_0_0_9), .A1 (n_0_0_12), .A2 (n_0_0_10), .B1 (\values[9] [15] ), .B2 (n_0_0_63));
INV_X1 i_0_0_13 (.ZN (n_0_0_8), .A (n_0_0_9));
AOI21_X1 i_0_0_12 (.ZN (n_0_0_7), .A (n_0_0_9), .B1 (n_0_0_65), .B2 (n_0_0_66));
INV_X2 i_0_0_11 (.ZN (n_0_0_6), .A (n_0_0_7));
NOR2_X4 i_0_0_10 (.ZN (spt__n4), .A1 (n_0_0_118), .A2 (n_0_0_6));
NAND2_X1 i_0_0_9 (.ZN (class_out[3]), .A1 (n_0_0_7), .A2 (n_0_0_118));
AOI21_X1 i_0_0_8 (.ZN (class_out[2]), .A (n_0_0_6), .B1 (n_0_0_119), .B2 (n_0_0_345));
OAI21_X1 i_0_0_7 (.ZN (n_0_0_5), .A (n_0_0_237), .B1 (n_0_0_347), .B2 (n_0_0_354));
AOI21_X1 i_0_0_6 (.ZN (class_out[1]), .A (n_0_0_6), .B1 (n_0_0_5), .B2 (n_0_0_120));
OAI21_X1 i_0_0_5 (.ZN (n_0_0_4), .A (spw__n671), .B1 (n_0_0_349), .B2 (n_0_0_479));
AOI21_X1 i_0_0_4 (.ZN (n_0_0_3), .A (n_0_0_292), .B1 (n_0_0_4), .B2 (spw__n698));
OAI21_X1 i_0_0_3 (.ZN (n_0_0_2), .A (n_0_0_178), .B1 (n_0_0_3), .B2 (n_0_0_238));
INV_X1 i_0_0_2 (.ZN (n_0_0_1), .A (n_0_0_2));
OAI21_X1 i_0_0_1 (.ZN (n_0_0_0), .A (n_0_0_64), .B1 (n_0_0_1), .B2 (n_0_0_121));
NAND2_X1 i_0_0_0 (.ZN (class_out[0]), .A1 (n_0_0_8), .A2 (n_0_0_0));
BUF_X4 spt__c1 (.Z (n_0_0_64), .A (spt__n1));
BUF_X4 spt__c4 (.Z (class_out[4]), .A (spt__n4));
BUF_X4 spt__c7 (.Z (n_0_0_121), .A (spt__n7));
BUF_X4 spw__c46 (.Z (n_0_0_479), .A (spw__n46));
BUF_X1 spw__L1_c642 (.Z (spw__n644), .A (n_0_0_478));
BUF_X2 spw__L2_c643 (.Z (spw__n645), .A (spw__n644));
BUF_X2 spw__L3_c644 (.Z (spw__n646), .A (spw__n645));
BUF_X1 spw__L1_c669 (.Z (spw__n671), .A (n_0_0_417));
BUF_X2 spw__L2_c670 (.Z (spw__n672), .A (spw__n671));
BUF_X1 spw__L1_c696 (.Z (spw__n698), .A (n_0_0_355));
BUF_X2 spw__c683 (.Z (n_0_0_402), .A (spw__n685));

endmodule //Softmax


