/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sun May 23 15:17:31 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1797485097 */

module datapath__0_120(mem_idx, p_0);
   input [31:0]mem_idx;
   output [31:0]p_0;

   HA_X1 i_0 (.A(mem_idx[1]), .B(mem_idx[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(mem_idx[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_2 (.A(mem_idx[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_3 (.A(mem_idx[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_4 (.A(mem_idx[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_5 (.A(mem_idx[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_6 (.A(mem_idx[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_7 (.A(mem_idx[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_8 (.A(mem_idx[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_9 (.A(mem_idx[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_10 (.A(mem_idx[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_11 (.A(mem_idx[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_12 (.A(mem_idx[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_13 (.A(mem_idx[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_14 (.A(mem_idx[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_15 (.A(mem_idx[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_16 (.A(mem_idx[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_17 (.A(mem_idx[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_18 (.A(mem_idx[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_19 (.A(mem_idx[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_20 (.A(mem_idx[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_21 (.A(mem_idx[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_22 (.A(mem_idx[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_23 (.A(mem_idx[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_24 (.A(mem_idx[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_25 (.A(mem_idx[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_26 (.A(mem_idx[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_27 (.A(mem_idx[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_28 (.A(mem_idx[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_29 (.A(mem_idx[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_30 (.A(mem_idx[31]), .B(n_29), .Z(p_0[31]));
endmodule

module DMA(i_read, i_address, i_count, clk, i_mem_data, o_mem_addr, 
      \o_buffer[119] , \o_buffer[118] , \o_buffer[117] , \o_buffer[116] , 
      \o_buffer[115] , \o_buffer[114] , \o_buffer[113] , \o_buffer[112] , 
      \o_buffer[111] , \o_buffer[110] , \o_buffer[109] , \o_buffer[108] , 
      \o_buffer[107] , \o_buffer[106] , \o_buffer[105] , \o_buffer[104] , 
      \o_buffer[103] , \o_buffer[102] , \o_buffer[101] , \o_buffer[100] , 
      \o_buffer[99] , \o_buffer[98] , \o_buffer[97] , \o_buffer[96] , 
      \o_buffer[95] , \o_buffer[94] , \o_buffer[93] , \o_buffer[92] , 
      \o_buffer[91] , \o_buffer[90] , \o_buffer[89] , \o_buffer[88] , 
      \o_buffer[87] , \o_buffer[86] , \o_buffer[85] , \o_buffer[84] , 
      \o_buffer[83] , \o_buffer[82] , \o_buffer[81] , \o_buffer[80] , 
      \o_buffer[79] , \o_buffer[78] , \o_buffer[77] , \o_buffer[76] , 
      \o_buffer[75] , \o_buffer[74] , \o_buffer[73] , \o_buffer[72] , 
      \o_buffer[71] , \o_buffer[70] , \o_buffer[69] , \o_buffer[68] , 
      \o_buffer[67] , \o_buffer[66] , \o_buffer[65] , \o_buffer[64] , 
      \o_buffer[63] , \o_buffer[62] , \o_buffer[61] , \o_buffer[60] , 
      \o_buffer[59] , \o_buffer[58] , \o_buffer[57] , \o_buffer[56] , 
      \o_buffer[55] , \o_buffer[54] , \o_buffer[53] , \o_buffer[52] , 
      \o_buffer[51] , \o_buffer[50] , \o_buffer[49] , \o_buffer[48] , 
      \o_buffer[47] , \o_buffer[46] , \o_buffer[45] , \o_buffer[44] , 
      \o_buffer[43] , \o_buffer[42] , \o_buffer[41] , \o_buffer[40] , 
      \o_buffer[39] , \o_buffer[38] , \o_buffer[37] , \o_buffer[36] , 
      \o_buffer[35] , \o_buffer[34] , \o_buffer[33] , \o_buffer[32] , 
      \o_buffer[31] , \o_buffer[30] , \o_buffer[29] , \o_buffer[28] , 
      \o_buffer[27] , \o_buffer[26] , \o_buffer[25] , \o_buffer[24] , 
      \o_buffer[23] , \o_buffer[22] , \o_buffer[21] , \o_buffer[20] , 
      \o_buffer[19] , \o_buffer[18] , \o_buffer[17] , \o_buffer[16] , 
      \o_buffer[15] , \o_buffer[14] , \o_buffer[13] , \o_buffer[12] , 
      \o_buffer[11] , \o_buffer[10] , \o_buffer[9] , \o_buffer[8] , 
      \o_buffer[7] , \o_buffer[6] , \o_buffer[5] , \o_buffer[4] , \o_buffer[3] , 
      \o_buffer[2] , \o_buffer[1] , \o_buffer[0] , o_ready);
   input i_read;
   input [9:0]i_address;
   input [9:0]i_count;
   input clk;
   input [15:0]i_mem_data;
   output [9:0]o_mem_addr;
   output [15:0]\o_buffer[119] ;
   output [15:0]\o_buffer[118] ;
   output [15:0]\o_buffer[117] ;
   output [15:0]\o_buffer[116] ;
   output [15:0]\o_buffer[115] ;
   output [15:0]\o_buffer[114] ;
   output [15:0]\o_buffer[113] ;
   output [15:0]\o_buffer[112] ;
   output [15:0]\o_buffer[111] ;
   output [15:0]\o_buffer[110] ;
   output [15:0]\o_buffer[109] ;
   output [15:0]\o_buffer[108] ;
   output [15:0]\o_buffer[107] ;
   output [15:0]\o_buffer[106] ;
   output [15:0]\o_buffer[105] ;
   output [15:0]\o_buffer[104] ;
   output [15:0]\o_buffer[103] ;
   output [15:0]\o_buffer[102] ;
   output [15:0]\o_buffer[101] ;
   output [15:0]\o_buffer[100] ;
   output [15:0]\o_buffer[99] ;
   output [15:0]\o_buffer[98] ;
   output [15:0]\o_buffer[97] ;
   output [15:0]\o_buffer[96] ;
   output [15:0]\o_buffer[95] ;
   output [15:0]\o_buffer[94] ;
   output [15:0]\o_buffer[93] ;
   output [15:0]\o_buffer[92] ;
   output [15:0]\o_buffer[91] ;
   output [15:0]\o_buffer[90] ;
   output [15:0]\o_buffer[89] ;
   output [15:0]\o_buffer[88] ;
   output [15:0]\o_buffer[87] ;
   output [15:0]\o_buffer[86] ;
   output [15:0]\o_buffer[85] ;
   output [15:0]\o_buffer[84] ;
   output [15:0]\o_buffer[83] ;
   output [15:0]\o_buffer[82] ;
   output [15:0]\o_buffer[81] ;
   output [15:0]\o_buffer[80] ;
   output [15:0]\o_buffer[79] ;
   output [15:0]\o_buffer[78] ;
   output [15:0]\o_buffer[77] ;
   output [15:0]\o_buffer[76] ;
   output [15:0]\o_buffer[75] ;
   output [15:0]\o_buffer[74] ;
   output [15:0]\o_buffer[73] ;
   output [15:0]\o_buffer[72] ;
   output [15:0]\o_buffer[71] ;
   output [15:0]\o_buffer[70] ;
   output [15:0]\o_buffer[69] ;
   output [15:0]\o_buffer[68] ;
   output [15:0]\o_buffer[67] ;
   output [15:0]\o_buffer[66] ;
   output [15:0]\o_buffer[65] ;
   output [15:0]\o_buffer[64] ;
   output [15:0]\o_buffer[63] ;
   output [15:0]\o_buffer[62] ;
   output [15:0]\o_buffer[61] ;
   output [15:0]\o_buffer[60] ;
   output [15:0]\o_buffer[59] ;
   output [15:0]\o_buffer[58] ;
   output [15:0]\o_buffer[57] ;
   output [15:0]\o_buffer[56] ;
   output [15:0]\o_buffer[55] ;
   output [15:0]\o_buffer[54] ;
   output [15:0]\o_buffer[53] ;
   output [15:0]\o_buffer[52] ;
   output [15:0]\o_buffer[51] ;
   output [15:0]\o_buffer[50] ;
   output [15:0]\o_buffer[49] ;
   output [15:0]\o_buffer[48] ;
   output [15:0]\o_buffer[47] ;
   output [15:0]\o_buffer[46] ;
   output [15:0]\o_buffer[45] ;
   output [15:0]\o_buffer[44] ;
   output [15:0]\o_buffer[43] ;
   output [15:0]\o_buffer[42] ;
   output [15:0]\o_buffer[41] ;
   output [15:0]\o_buffer[40] ;
   output [15:0]\o_buffer[39] ;
   output [15:0]\o_buffer[38] ;
   output [15:0]\o_buffer[37] ;
   output [15:0]\o_buffer[36] ;
   output [15:0]\o_buffer[35] ;
   output [15:0]\o_buffer[34] ;
   output [15:0]\o_buffer[33] ;
   output [15:0]\o_buffer[32] ;
   output [15:0]\o_buffer[31] ;
   output [15:0]\o_buffer[30] ;
   output [15:0]\o_buffer[29] ;
   output [15:0]\o_buffer[28] ;
   output [15:0]\o_buffer[27] ;
   output [15:0]\o_buffer[26] ;
   output [15:0]\o_buffer[25] ;
   output [15:0]\o_buffer[24] ;
   output [15:0]\o_buffer[23] ;
   output [15:0]\o_buffer[22] ;
   output [15:0]\o_buffer[21] ;
   output [15:0]\o_buffer[20] ;
   output [15:0]\o_buffer[19] ;
   output [15:0]\o_buffer[18] ;
   output [15:0]\o_buffer[17] ;
   output [15:0]\o_buffer[16] ;
   output [15:0]\o_buffer[15] ;
   output [15:0]\o_buffer[14] ;
   output [15:0]\o_buffer[13] ;
   output [15:0]\o_buffer[12] ;
   output [15:0]\o_buffer[11] ;
   output [15:0]\o_buffer[10] ;
   output [15:0]\o_buffer[9] ;
   output [15:0]\o_buffer[8] ;
   output [15:0]\o_buffer[7] ;
   output [15:0]\o_buffer[6] ;
   output [15:0]\o_buffer[5] ;
   output [15:0]\o_buffer[4] ;
   output [15:0]\o_buffer[3] ;
   output [15:0]\o_buffer[2] ;
   output [15:0]\o_buffer[1] ;
   output [15:0]\o_buffer[0] ;
   output o_ready;

   wire n_123_959;
   wire n_123_958;
   wire n_123_957;
   wire n_123_956;
   wire n_123_955;
   wire n_123_954;
   wire n_123_953;
   wire n_123_952;
   wire n_123_951;
   wire n_123_950;
   wire n_123_949;
   wire n_123_948;
   wire n_123_947;
   wire n_123_946;
   wire n_123_945;
   wire n_123_944;
   wire n_123_943;
   wire n_123_942;
   wire n_123_941;
   wire n_123_940;
   wire n_123_939;
   wire n_123_938;
   wire n_123_937;
   wire n_123_936;
   wire n_123_935;
   wire n_123_934;
   wire n_123_933;
   wire n_123_932;
   wire n_123_931;
   wire n_123_930;
   wire n_123_929;
   wire n_123_928;
   wire n_123_927;
   wire n_123_926;
   wire n_123_925;
   wire n_123_924;
   wire n_123_923;
   wire n_123_922;
   wire n_123_921;
   wire n_123_920;
   wire n_123_919;
   wire n_123_918;
   wire n_123_917;
   wire n_123_916;
   wire n_123_915;
   wire n_123_914;
   wire n_123_913;
   wire n_123_912;
   wire n_123_911;
   wire n_123_910;
   wire n_123_909;
   wire n_123_908;
   wire n_123_907;
   wire n_123_906;
   wire n_123_905;
   wire n_123_904;
   wire n_123_903;
   wire n_123_902;
   wire n_123_901;
   wire n_123_900;
   wire n_123_899;
   wire n_123_898;
   wire n_123_897;
   wire n_123_896;
   wire n_123_895;
   wire n_123_894;
   wire n_123_893;
   wire n_123_892;
   wire n_123_891;
   wire n_123_890;
   wire n_123_889;
   wire n_123_888;
   wire n_123_887;
   wire n_123_886;
   wire n_123_885;
   wire n_123_884;
   wire n_123_883;
   wire n_123_882;
   wire n_123_881;
   wire n_123_880;
   wire n_123_879;
   wire n_123_878;
   wire n_123_877;
   wire n_123_876;
   wire n_123_875;
   wire n_123_874;
   wire n_123_873;
   wire n_123_872;
   wire n_123_871;
   wire n_123_870;
   wire n_123_869;
   wire n_123_868;
   wire n_123_867;
   wire n_123_866;
   wire n_123_865;
   wire n_123_864;
   wire n_123_863;
   wire n_123_862;
   wire n_123_861;
   wire n_123_860;
   wire n_123_859;
   wire n_123_858;
   wire n_123_857;
   wire n_123_856;
   wire n_123_855;
   wire n_123_854;
   wire n_123_853;
   wire n_123_852;
   wire n_123_851;
   wire n_123_850;
   wire n_123_849;
   wire n_123_848;
   wire n_123_847;
   wire n_123_846;
   wire n_123_845;
   wire n_123_844;
   wire n_123_843;
   wire n_123_842;
   wire n_123_841;
   wire n_123_840;
   wire n_123_839;
   wire n_123_838;
   wire n_123_837;
   wire n_123_836;
   wire n_123_835;
   wire n_123_834;
   wire n_123_833;
   wire n_123_832;
   wire n_123_831;
   wire n_123_830;
   wire n_123_829;
   wire n_123_828;
   wire n_123_827;
   wire n_123_826;
   wire n_123_825;
   wire n_123_824;
   wire n_123_823;
   wire n_123_822;
   wire n_123_821;
   wire n_123_820;
   wire n_123_819;
   wire n_123_818;
   wire n_123_817;
   wire n_123_816;
   wire n_123_815;
   wire n_123_814;
   wire n_123_813;
   wire n_123_812;
   wire n_123_811;
   wire n_123_810;
   wire n_123_809;
   wire n_123_808;
   wire n_123_807;
   wire n_123_806;
   wire n_123_805;
   wire n_123_804;
   wire n_123_803;
   wire n_123_802;
   wire n_123_801;
   wire n_123_800;
   wire n_123_799;
   wire n_123_798;
   wire n_123_797;
   wire n_123_796;
   wire n_123_795;
   wire n_123_794;
   wire n_123_793;
   wire n_123_792;
   wire n_123_791;
   wire n_123_790;
   wire n_123_789;
   wire n_123_788;
   wire n_123_787;
   wire n_123_786;
   wire n_123_785;
   wire n_123_784;
   wire n_123_783;
   wire n_123_782;
   wire n_123_781;
   wire n_123_780;
   wire n_123_779;
   wire n_123_778;
   wire n_123_777;
   wire n_123_776;
   wire n_123_775;
   wire n_123_774;
   wire n_123_773;
   wire n_123_772;
   wire n_123_771;
   wire n_123_770;
   wire n_123_769;
   wire n_123_768;
   wire n_123_767;
   wire n_123_766;
   wire n_123_765;
   wire n_123_764;
   wire n_123_763;
   wire n_123_762;
   wire n_123_761;
   wire n_123_760;
   wire n_123_759;
   wire n_123_758;
   wire n_123_757;
   wire n_123_756;
   wire n_123_755;
   wire n_123_754;
   wire n_123_753;
   wire n_123_752;
   wire n_123_751;
   wire n_123_750;
   wire n_123_749;
   wire n_123_748;
   wire n_123_747;
   wire n_123_746;
   wire n_123_745;
   wire n_123_744;
   wire n_123_743;
   wire n_123_742;
   wire n_123_741;
   wire n_123_740;
   wire n_123_739;
   wire n_123_738;
   wire n_123_737;
   wire n_123_736;
   wire n_123_735;
   wire n_123_734;
   wire n_123_733;
   wire n_123_732;
   wire n_123_731;
   wire n_123_730;
   wire n_123_729;
   wire n_123_728;
   wire n_123_727;
   wire n_123_726;
   wire n_123_725;
   wire n_123_724;
   wire n_123_723;
   wire n_123_722;
   wire n_123_721;
   wire n_123_720;
   wire n_123_719;
   wire n_123_718;
   wire n_123_717;
   wire n_123_716;
   wire n_123_715;
   wire n_123_714;
   wire n_123_713;
   wire n_123_712;
   wire n_123_711;
   wire n_123_710;
   wire n_123_709;
   wire n_123_708;
   wire n_123_707;
   wire n_123_706;
   wire n_123_705;
   wire n_123_704;
   wire n_123_703;
   wire n_123_702;
   wire n_123_701;
   wire n_123_700;
   wire n_123_699;
   wire n_123_698;
   wire n_123_697;
   wire n_123_696;
   wire n_123_695;
   wire n_123_694;
   wire n_123_693;
   wire n_123_692;
   wire n_123_691;
   wire n_123_690;
   wire n_123_689;
   wire n_123_688;
   wire n_123_687;
   wire n_123_686;
   wire n_123_685;
   wire n_123_684;
   wire n_123_683;
   wire n_123_682;
   wire n_123_681;
   wire n_123_680;
   wire n_123_679;
   wire n_123_678;
   wire n_123_677;
   wire n_123_676;
   wire n_123_675;
   wire n_123_674;
   wire n_123_673;
   wire n_123_672;
   wire n_123_671;
   wire n_123_670;
   wire n_123_669;
   wire n_123_668;
   wire n_123_667;
   wire n_123_666;
   wire n_123_665;
   wire n_123_664;
   wire n_123_663;
   wire n_123_662;
   wire n_123_661;
   wire n_123_660;
   wire n_123_659;
   wire n_123_658;
   wire n_123_657;
   wire n_123_656;
   wire n_123_655;
   wire n_123_654;
   wire n_123_653;
   wire n_123_652;
   wire n_123_651;
   wire n_123_650;
   wire n_123_649;
   wire n_123_648;
   wire n_123_647;
   wire n_123_646;
   wire n_123_645;
   wire n_123_644;
   wire n_123_643;
   wire n_123_642;
   wire n_123_641;
   wire n_123_640;
   wire n_123_639;
   wire n_123_638;
   wire n_123_637;
   wire n_123_636;
   wire n_123_635;
   wire n_123_634;
   wire n_123_633;
   wire n_123_632;
   wire n_123_631;
   wire n_123_630;
   wire n_123_629;
   wire n_123_628;
   wire n_123_627;
   wire n_123_626;
   wire n_123_625;
   wire n_123_624;
   wire n_123_623;
   wire n_123_622;
   wire n_123_621;
   wire n_123_620;
   wire n_123_619;
   wire n_123_618;
   wire n_123_617;
   wire n_123_616;
   wire n_123_615;
   wire n_123_614;
   wire n_123_613;
   wire n_123_612;
   wire n_123_611;
   wire n_123_610;
   wire n_123_609;
   wire n_123_608;
   wire n_123_607;
   wire n_123_606;
   wire n_123_605;
   wire n_123_604;
   wire n_123_603;
   wire n_123_602;
   wire n_123_601;
   wire n_123_600;
   wire n_123_599;
   wire n_123_598;
   wire n_123_597;
   wire n_123_596;
   wire n_123_595;
   wire n_123_594;
   wire n_123_593;
   wire n_123_592;
   wire n_123_591;
   wire n_123_590;
   wire n_123_589;
   wire n_123_588;
   wire n_123_587;
   wire n_123_586;
   wire n_123_585;
   wire n_123_584;
   wire n_123_583;
   wire n_123_582;
   wire n_123_581;
   wire n_123_580;
   wire n_123_579;
   wire n_123_578;
   wire n_123_577;
   wire n_123_576;
   wire n_123_575;
   wire n_123_574;
   wire n_123_573;
   wire n_123_572;
   wire n_123_571;
   wire n_123_570;
   wire n_123_569;
   wire n_123_568;
   wire n_123_567;
   wire n_123_566;
   wire n_123_565;
   wire n_123_564;
   wire n_123_563;
   wire n_123_562;
   wire n_123_561;
   wire n_123_560;
   wire n_123_559;
   wire n_123_558;
   wire n_123_557;
   wire n_123_556;
   wire n_123_555;
   wire n_123_554;
   wire n_123_553;
   wire n_123_552;
   wire n_123_551;
   wire n_123_550;
   wire n_123_549;
   wire n_123_548;
   wire n_123_547;
   wire n_123_546;
   wire n_123_545;
   wire n_123_544;
   wire n_123_543;
   wire n_123_542;
   wire n_123_541;
   wire n_123_540;
   wire n_123_539;
   wire n_123_538;
   wire n_123_537;
   wire n_123_536;
   wire n_123_535;
   wire n_123_534;
   wire n_123_533;
   wire n_123_532;
   wire n_123_531;
   wire n_123_530;
   wire n_123_529;
   wire n_123_528;
   wire n_123_527;
   wire n_123_526;
   wire n_123_525;
   wire n_123_524;
   wire n_123_523;
   wire n_123_522;
   wire n_123_521;
   wire n_123_520;
   wire n_123_519;
   wire n_123_518;
   wire n_123_517;
   wire n_123_516;
   wire n_123_515;
   wire n_123_514;
   wire n_123_513;
   wire n_123_512;
   wire n_123_511;
   wire n_123_510;
   wire n_123_509;
   wire n_123_508;
   wire n_123_507;
   wire n_123_506;
   wire n_123_505;
   wire n_123_504;
   wire n_123_503;
   wire n_123_502;
   wire n_123_501;
   wire n_123_500;
   wire n_123_499;
   wire n_123_498;
   wire n_123_497;
   wire n_123_496;
   wire n_123_495;
   wire n_123_494;
   wire n_123_493;
   wire n_123_492;
   wire n_123_491;
   wire n_123_490;
   wire n_123_489;
   wire n_123_488;
   wire n_123_487;
   wire n_123_486;
   wire n_123_485;
   wire n_123_484;
   wire n_123_483;
   wire n_123_482;
   wire n_123_481;
   wire n_123_480;
   wire n_123_479;
   wire n_123_478;
   wire n_123_477;
   wire n_123_476;
   wire n_123_475;
   wire n_123_474;
   wire n_123_473;
   wire n_123_472;
   wire n_123_471;
   wire n_123_470;
   wire n_123_469;
   wire n_123_468;
   wire n_123_467;
   wire n_123_466;
   wire n_123_465;
   wire n_123_464;
   wire n_123_463;
   wire n_123_462;
   wire n_123_461;
   wire n_123_460;
   wire n_123_459;
   wire n_123_458;
   wire n_123_457;
   wire n_123_456;
   wire n_123_455;
   wire n_123_454;
   wire n_123_453;
   wire n_123_452;
   wire n_123_451;
   wire n_123_450;
   wire n_123_449;
   wire n_123_448;
   wire n_123_447;
   wire n_123_446;
   wire n_123_445;
   wire n_123_444;
   wire n_123_443;
   wire n_123_442;
   wire n_123_441;
   wire n_123_440;
   wire n_123_439;
   wire n_123_438;
   wire n_123_437;
   wire n_123_436;
   wire n_123_435;
   wire n_123_434;
   wire n_123_433;
   wire n_123_432;
   wire n_123_431;
   wire n_123_430;
   wire n_123_429;
   wire n_123_428;
   wire n_123_427;
   wire n_123_426;
   wire n_123_425;
   wire n_123_424;
   wire n_123_423;
   wire n_123_422;
   wire n_123_421;
   wire n_123_420;
   wire n_123_419;
   wire n_123_418;
   wire n_123_417;
   wire n_123_416;
   wire n_123_415;
   wire n_123_414;
   wire n_123_413;
   wire n_123_412;
   wire n_123_411;
   wire n_123_410;
   wire n_123_409;
   wire n_123_408;
   wire n_123_407;
   wire n_123_406;
   wire n_123_405;
   wire n_123_404;
   wire n_123_403;
   wire n_123_402;
   wire n_123_401;
   wire n_123_400;
   wire n_123_399;
   wire n_123_398;
   wire n_123_397;
   wire n_123_396;
   wire n_123_395;
   wire n_123_394;
   wire n_123_393;
   wire n_123_392;
   wire n_123_391;
   wire n_123_390;
   wire n_123_389;
   wire n_123_388;
   wire n_123_387;
   wire n_123_386;
   wire n_123_385;
   wire n_123_384;
   wire n_123_383;
   wire n_123_382;
   wire n_123_381;
   wire n_123_380;
   wire n_123_379;
   wire n_123_378;
   wire n_123_377;
   wire n_123_376;
   wire n_123_375;
   wire n_123_374;
   wire n_123_373;
   wire n_123_372;
   wire n_123_371;
   wire n_123_370;
   wire n_123_369;
   wire n_123_368;
   wire n_123_367;
   wire n_123_366;
   wire n_123_365;
   wire n_123_364;
   wire n_123_363;
   wire n_123_362;
   wire n_123_361;
   wire n_123_360;
   wire n_123_359;
   wire n_123_358;
   wire n_123_357;
   wire n_123_356;
   wire n_123_355;
   wire n_123_354;
   wire n_123_353;
   wire n_123_352;
   wire n_123_351;
   wire n_123_350;
   wire n_123_349;
   wire n_123_348;
   wire n_123_347;
   wire n_123_346;
   wire n_123_345;
   wire n_123_344;
   wire n_123_343;
   wire n_123_342;
   wire n_123_341;
   wire n_123_340;
   wire n_123_339;
   wire n_123_338;
   wire n_123_337;
   wire n_123_336;
   wire n_123_335;
   wire n_123_334;
   wire n_123_333;
   wire n_123_332;
   wire n_123_331;
   wire n_123_330;
   wire n_123_329;
   wire n_123_328;
   wire n_123_327;
   wire n_123_326;
   wire n_123_325;
   wire n_123_324;
   wire n_123_323;
   wire n_123_322;
   wire n_123_321;
   wire n_123_320;
   wire n_123_319;
   wire n_123_318;
   wire n_123_317;
   wire n_123_316;
   wire n_123_315;
   wire n_123_314;
   wire n_123_313;
   wire n_123_312;
   wire n_123_311;
   wire n_123_310;
   wire n_123_309;
   wire n_123_308;
   wire n_123_307;
   wire n_123_306;
   wire n_123_305;
   wire n_123_304;
   wire n_123_303;
   wire n_123_302;
   wire n_123_301;
   wire n_123_300;
   wire n_123_299;
   wire n_123_298;
   wire n_123_297;
   wire n_123_296;
   wire n_123_295;
   wire n_123_294;
   wire n_123_293;
   wire n_123_292;
   wire n_123_291;
   wire n_123_290;
   wire n_123_289;
   wire n_123_288;
   wire n_123_287;
   wire n_123_286;
   wire n_123_285;
   wire n_123_284;
   wire n_123_283;
   wire n_123_282;
   wire n_123_281;
   wire n_123_280;
   wire n_123_279;
   wire n_123_278;
   wire n_123_277;
   wire n_123_276;
   wire n_123_275;
   wire n_123_274;
   wire n_123_273;
   wire n_123_272;
   wire n_123_271;
   wire n_123_270;
   wire n_123_269;
   wire n_123_268;
   wire n_123_267;
   wire n_123_266;
   wire n_123_265;
   wire n_123_264;
   wire n_123_263;
   wire n_123_262;
   wire n_123_261;
   wire n_123_260;
   wire n_123_259;
   wire n_123_258;
   wire n_123_257;
   wire n_123_256;
   wire n_123_255;
   wire n_123_254;
   wire n_123_253;
   wire n_123_252;
   wire n_123_251;
   wire n_123_250;
   wire n_123_249;
   wire n_123_248;
   wire n_123_247;
   wire n_123_246;
   wire n_123_245;
   wire n_123_244;
   wire n_123_243;
   wire n_123_242;
   wire n_123_241;
   wire n_123_240;
   wire n_123_239;
   wire n_123_238;
   wire n_123_237;
   wire n_123_236;
   wire n_123_235;
   wire n_123_234;
   wire n_123_233;
   wire n_123_232;
   wire n_123_231;
   wire n_123_230;
   wire n_123_229;
   wire n_123_228;
   wire n_123_227;
   wire n_123_226;
   wire n_123_225;
   wire n_123_224;
   wire n_123_223;
   wire n_123_222;
   wire n_123_221;
   wire n_123_220;
   wire n_123_219;
   wire n_123_218;
   wire n_123_217;
   wire n_123_216;
   wire n_123_215;
   wire n_123_214;
   wire n_123_213;
   wire n_123_212;
   wire n_123_211;
   wire n_123_210;
   wire n_123_209;
   wire n_123_208;
   wire n_123_207;
   wire n_123_206;
   wire n_123_205;
   wire n_123_204;
   wire n_123_203;
   wire n_123_202;
   wire n_123_201;
   wire n_123_200;
   wire n_123_199;
   wire n_123_198;
   wire n_123_197;
   wire n_123_196;
   wire n_123_195;
   wire n_123_194;
   wire n_123_193;
   wire n_123_192;
   wire n_123_191;
   wire n_123_190;
   wire n_123_189;
   wire n_123_188;
   wire n_123_187;
   wire n_123_186;
   wire n_123_185;
   wire n_123_184;
   wire n_123_183;
   wire n_123_182;
   wire n_123_181;
   wire n_123_180;
   wire n_123_179;
   wire n_123_178;
   wire n_123_177;
   wire n_123_176;
   wire n_123_175;
   wire n_123_174;
   wire n_123_173;
   wire n_123_172;
   wire n_123_171;
   wire n_123_170;
   wire n_123_169;
   wire n_123_168;
   wire n_123_167;
   wire n_123_166;
   wire n_123_165;
   wire n_123_164;
   wire n_123_163;
   wire n_123_162;
   wire n_123_161;
   wire n_123_160;
   wire n_123_159;
   wire n_123_158;
   wire n_123_157;
   wire n_123_156;
   wire n_123_155;
   wire n_123_154;
   wire n_123_153;
   wire n_123_152;
   wire n_123_151;
   wire n_123_150;
   wire n_123_149;
   wire n_123_148;
   wire n_123_147;
   wire n_123_146;
   wire n_123_145;
   wire n_123_144;
   wire n_123_143;
   wire n_123_142;
   wire n_123_141;
   wire n_123_140;
   wire n_123_139;
   wire n_123_138;
   wire n_123_137;
   wire n_123_136;
   wire n_123_135;
   wire n_123_134;
   wire n_123_133;
   wire n_123_132;
   wire n_123_131;
   wire n_123_130;
   wire n_123_129;
   wire n_123_128;
   wire n_123_127;
   wire n_123_126;
   wire n_123_125;
   wire n_123_124;
   wire n_123_123;
   wire n_123_122;
   wire n_123_121;
   wire n_123_120;
   wire n_123_119;
   wire n_123_118;
   wire n_123_117;
   wire n_123_116;
   wire n_123_115;
   wire n_123_114;
   wire n_123_113;
   wire n_123_112;
   wire n_123_111;
   wire n_123_110;
   wire n_123_109;
   wire n_123_108;
   wire n_123_107;
   wire n_123_106;
   wire n_123_105;
   wire n_123_104;
   wire n_123_103;
   wire n_123_102;
   wire n_123_101;
   wire n_123_100;
   wire n_123_99;
   wire n_123_98;
   wire n_123_97;
   wire n_123_96;
   wire n_123_95;
   wire n_123_94;
   wire n_123_93;
   wire n_123_92;
   wire n_123_91;
   wire n_123_90;
   wire n_123_89;
   wire n_123_88;
   wire n_123_87;
   wire n_123_86;
   wire n_123_85;
   wire n_123_84;
   wire n_123_83;
   wire n_123_82;
   wire n_123_81;
   wire n_123_80;
   wire n_123_79;
   wire n_123_78;
   wire n_123_77;
   wire n_123_76;
   wire n_123_75;
   wire n_123_74;
   wire n_123_73;
   wire n_123_72;
   wire n_123_71;
   wire n_123_70;
   wire n_123_69;
   wire n_123_68;
   wire n_123_67;
   wire n_123_66;
   wire n_123_65;
   wire n_123_64;
   wire n_123_63;
   wire n_123_62;
   wire n_123_61;
   wire n_123_60;
   wire n_123_59;
   wire n_123_58;
   wire n_123_57;
   wire n_123_56;
   wire n_123_55;
   wire n_123_54;
   wire n_123_53;
   wire n_123_52;
   wire n_123_51;
   wire n_123_50;
   wire n_123_49;
   wire n_123_48;
   wire n_123_47;
   wire n_123_46;
   wire n_123_45;
   wire n_123_44;
   wire n_123_43;
   wire n_123_42;
   wire n_123_41;
   wire n_123_40;
   wire n_123_39;
   wire n_123_38;
   wire n_123_37;
   wire n_123_36;
   wire n_123_35;
   wire n_123_34;
   wire n_123_33;
   wire n_123_32;
   wire n_123_31;
   wire n_123_30;
   wire n_123_29;
   wire n_123_28;
   wire n_123_27;
   wire n_123_26;
   wire n_123_25;
   wire n_123_24;
   wire n_123_23;
   wire n_123_22;
   wire n_123_21;
   wire n_123_20;
   wire n_123_19;
   wire n_123_18;
   wire n_123_17;
   wire n_123_16;
   wire n_123_15;
   wire n_123_14;
   wire n_123_13;
   wire n_123_12;
   wire n_123_11;
   wire n_123_10;
   wire n_123_9;
   wire n_123_8;
   wire n_123_7;
   wire n_123_6;
   wire n_123_5;
   wire n_123_4;
   wire n_123_3;
   wire n_123_2;
   wire n_123_1;
   wire n_123_0;
   wire n_132_959;
   wire n_132_958;
   wire n_132_957;
   wire n_132_956;
   wire n_132_955;
   wire n_132_954;
   wire n_132_953;
   wire n_132_952;
   wire n_132_951;
   wire n_132_950;
   wire n_132_949;
   wire n_132_948;
   wire n_132_947;
   wire n_132_946;
   wire n_132_945;
   wire n_132_944;
   wire n_132_943;
   wire n_132_942;
   wire n_132_941;
   wire n_132_940;
   wire n_132_939;
   wire n_132_938;
   wire n_132_937;
   wire n_132_936;
   wire n_132_935;
   wire n_132_934;
   wire n_132_933;
   wire n_132_932;
   wire n_132_931;
   wire n_132_930;
   wire n_132_929;
   wire n_132_928;
   wire n_132_927;
   wire n_132_926;
   wire n_132_925;
   wire n_132_924;
   wire n_132_923;
   wire n_132_922;
   wire n_132_921;
   wire n_132_920;
   wire n_132_919;
   wire n_132_918;
   wire n_132_917;
   wire n_132_916;
   wire n_132_915;
   wire n_132_914;
   wire n_132_913;
   wire n_132_912;
   wire n_132_911;
   wire n_132_910;
   wire n_132_909;
   wire n_132_908;
   wire n_132_907;
   wire n_132_906;
   wire n_132_905;
   wire n_132_904;
   wire n_132_903;
   wire n_132_902;
   wire n_132_901;
   wire n_132_900;
   wire n_132_899;
   wire n_132_898;
   wire n_132_897;
   wire n_132_896;
   wire n_132_895;
   wire n_132_894;
   wire n_132_893;
   wire n_132_892;
   wire n_132_891;
   wire n_132_890;
   wire n_132_889;
   wire n_132_888;
   wire n_132_887;
   wire n_132_886;
   wire n_132_885;
   wire n_132_884;
   wire n_132_883;
   wire n_132_882;
   wire n_132_881;
   wire n_132_880;
   wire n_132_879;
   wire n_132_878;
   wire n_132_877;
   wire n_132_876;
   wire n_132_875;
   wire n_132_874;
   wire n_132_873;
   wire n_132_872;
   wire n_132_871;
   wire n_132_870;
   wire n_132_869;
   wire n_132_868;
   wire n_132_867;
   wire n_132_866;
   wire n_132_865;
   wire n_132_864;
   wire n_132_863;
   wire n_132_862;
   wire n_132_861;
   wire n_132_860;
   wire n_132_859;
   wire n_132_858;
   wire n_132_857;
   wire n_132_856;
   wire n_132_855;
   wire n_132_854;
   wire n_132_853;
   wire n_132_852;
   wire n_132_851;
   wire n_132_850;
   wire n_132_849;
   wire n_132_848;
   wire n_132_847;
   wire n_132_846;
   wire n_132_845;
   wire n_132_844;
   wire n_132_843;
   wire n_132_842;
   wire n_132_841;
   wire n_132_840;
   wire n_132_839;
   wire n_132_838;
   wire n_132_837;
   wire n_132_836;
   wire n_132_835;
   wire n_132_834;
   wire n_132_833;
   wire n_132_832;
   wire n_132_831;
   wire n_132_830;
   wire n_132_829;
   wire n_132_828;
   wire n_132_827;
   wire n_132_826;
   wire n_132_825;
   wire n_132_824;
   wire n_132_823;
   wire n_132_822;
   wire n_132_821;
   wire n_132_820;
   wire n_132_819;
   wire n_132_818;
   wire n_132_817;
   wire n_132_816;
   wire n_132_815;
   wire n_132_814;
   wire n_132_813;
   wire n_132_812;
   wire n_132_811;
   wire n_132_810;
   wire n_132_809;
   wire n_132_808;
   wire n_132_807;
   wire n_132_806;
   wire n_132_805;
   wire n_132_804;
   wire n_132_803;
   wire n_132_802;
   wire n_132_801;
   wire n_132_800;
   wire n_132_799;
   wire n_132_798;
   wire n_132_797;
   wire n_132_796;
   wire n_132_795;
   wire n_132_794;
   wire n_132_793;
   wire n_132_792;
   wire n_132_791;
   wire n_132_790;
   wire n_132_789;
   wire n_132_788;
   wire n_132_787;
   wire n_132_786;
   wire n_132_785;
   wire n_132_784;
   wire n_132_783;
   wire n_132_782;
   wire n_132_781;
   wire n_132_780;
   wire n_132_779;
   wire n_132_778;
   wire n_132_777;
   wire n_132_776;
   wire n_132_775;
   wire n_132_774;
   wire n_132_773;
   wire n_132_772;
   wire n_132_771;
   wire n_132_770;
   wire n_132_769;
   wire n_132_768;
   wire n_132_767;
   wire n_132_766;
   wire n_132_765;
   wire n_132_764;
   wire n_132_763;
   wire n_132_762;
   wire n_132_761;
   wire n_132_760;
   wire n_132_759;
   wire n_132_758;
   wire n_132_757;
   wire n_132_756;
   wire n_132_755;
   wire n_132_754;
   wire n_132_753;
   wire n_132_752;
   wire n_132_751;
   wire n_132_750;
   wire n_132_749;
   wire n_132_748;
   wire n_132_747;
   wire n_132_746;
   wire n_132_745;
   wire n_132_744;
   wire n_132_743;
   wire n_132_742;
   wire n_132_741;
   wire n_132_740;
   wire n_132_739;
   wire n_132_738;
   wire n_132_737;
   wire n_132_736;
   wire n_132_735;
   wire n_132_734;
   wire n_132_733;
   wire n_132_732;
   wire n_132_731;
   wire n_132_730;
   wire n_132_729;
   wire n_132_728;
   wire n_132_727;
   wire n_132_726;
   wire n_132_725;
   wire n_132_724;
   wire n_132_723;
   wire n_132_722;
   wire n_132_721;
   wire n_132_720;
   wire n_132_719;
   wire n_132_718;
   wire n_132_717;
   wire n_132_716;
   wire n_132_715;
   wire n_132_714;
   wire n_132_713;
   wire n_132_712;
   wire n_132_711;
   wire n_132_710;
   wire n_132_709;
   wire n_132_708;
   wire n_132_707;
   wire n_132_706;
   wire n_132_705;
   wire n_132_704;
   wire n_132_703;
   wire n_132_702;
   wire n_132_701;
   wire n_132_700;
   wire n_132_699;
   wire n_132_698;
   wire n_132_697;
   wire n_132_696;
   wire n_132_695;
   wire n_132_694;
   wire n_132_693;
   wire n_132_692;
   wire n_132_691;
   wire n_132_690;
   wire n_132_689;
   wire n_132_688;
   wire n_132_687;
   wire n_132_686;
   wire n_132_685;
   wire n_132_684;
   wire n_132_683;
   wire n_132_682;
   wire n_132_681;
   wire n_132_680;
   wire n_132_679;
   wire n_132_678;
   wire n_132_677;
   wire n_132_676;
   wire n_132_675;
   wire n_132_674;
   wire n_132_673;
   wire n_132_672;
   wire n_132_671;
   wire n_132_670;
   wire n_132_669;
   wire n_132_668;
   wire n_132_667;
   wire n_132_666;
   wire n_132_665;
   wire n_132_664;
   wire n_132_663;
   wire n_132_662;
   wire n_132_661;
   wire n_132_660;
   wire n_132_659;
   wire n_132_658;
   wire n_132_657;
   wire n_132_656;
   wire n_132_655;
   wire n_132_654;
   wire n_132_653;
   wire n_132_652;
   wire n_132_651;
   wire n_132_650;
   wire n_132_649;
   wire n_132_648;
   wire n_132_647;
   wire n_132_646;
   wire n_132_645;
   wire n_132_644;
   wire n_132_643;
   wire n_132_642;
   wire n_132_641;
   wire n_132_640;
   wire n_132_639;
   wire n_132_638;
   wire n_132_637;
   wire n_132_636;
   wire n_132_635;
   wire n_132_634;
   wire n_132_633;
   wire n_132_632;
   wire n_132_631;
   wire n_132_630;
   wire n_132_629;
   wire n_132_628;
   wire n_132_627;
   wire n_132_626;
   wire n_132_625;
   wire n_132_624;
   wire n_132_623;
   wire n_132_622;
   wire n_132_621;
   wire n_132_620;
   wire n_132_619;
   wire n_132_618;
   wire n_132_617;
   wire n_132_616;
   wire n_132_615;
   wire n_132_614;
   wire n_132_613;
   wire n_132_612;
   wire n_132_611;
   wire n_132_610;
   wire n_132_609;
   wire n_132_608;
   wire n_132_607;
   wire n_132_606;
   wire n_132_605;
   wire n_132_604;
   wire n_132_603;
   wire n_132_602;
   wire n_132_601;
   wire n_132_600;
   wire n_132_599;
   wire n_132_598;
   wire n_132_597;
   wire n_132_596;
   wire n_132_595;
   wire n_132_594;
   wire n_132_593;
   wire n_132_592;
   wire n_132_591;
   wire n_132_590;
   wire n_132_589;
   wire n_132_588;
   wire n_132_587;
   wire n_132_586;
   wire n_132_585;
   wire n_132_584;
   wire n_132_583;
   wire n_132_582;
   wire n_132_581;
   wire n_132_580;
   wire n_132_579;
   wire n_132_578;
   wire n_132_577;
   wire n_132_576;
   wire n_132_575;
   wire n_132_574;
   wire n_132_573;
   wire n_132_572;
   wire n_132_571;
   wire n_132_570;
   wire n_132_569;
   wire n_132_568;
   wire n_132_567;
   wire n_132_566;
   wire n_132_565;
   wire n_132_564;
   wire n_132_563;
   wire n_132_562;
   wire n_132_561;
   wire n_132_560;
   wire n_132_559;
   wire n_132_558;
   wire n_132_557;
   wire n_132_556;
   wire n_132_555;
   wire n_132_554;
   wire n_132_553;
   wire n_132_552;
   wire n_132_551;
   wire n_132_550;
   wire n_132_549;
   wire n_132_548;
   wire n_132_547;
   wire n_132_546;
   wire n_132_545;
   wire n_132_544;
   wire n_132_543;
   wire n_132_542;
   wire n_132_541;
   wire n_132_540;
   wire n_132_539;
   wire n_132_538;
   wire n_132_537;
   wire n_132_536;
   wire n_132_535;
   wire n_132_534;
   wire n_132_533;
   wire n_132_532;
   wire n_132_531;
   wire n_132_530;
   wire n_132_529;
   wire n_132_528;
   wire n_132_527;
   wire n_132_526;
   wire n_132_525;
   wire n_132_524;
   wire n_132_523;
   wire n_132_522;
   wire n_132_521;
   wire n_132_520;
   wire n_132_519;
   wire n_132_518;
   wire n_132_517;
   wire n_132_516;
   wire n_132_515;
   wire n_132_514;
   wire n_132_513;
   wire n_132_512;
   wire n_132_511;
   wire n_132_510;
   wire n_132_509;
   wire n_132_508;
   wire n_132_507;
   wire n_132_506;
   wire n_132_505;
   wire n_132_504;
   wire n_132_503;
   wire n_132_502;
   wire n_132_501;
   wire n_132_500;
   wire n_132_499;
   wire n_132_498;
   wire n_132_497;
   wire n_132_496;
   wire n_132_495;
   wire n_132_494;
   wire n_132_493;
   wire n_132_492;
   wire n_132_491;
   wire n_132_490;
   wire n_132_489;
   wire n_132_488;
   wire n_132_487;
   wire n_132_486;
   wire n_132_485;
   wire n_132_484;
   wire n_132_483;
   wire n_132_482;
   wire n_132_481;
   wire n_132_480;
   wire n_132_479;
   wire n_132_478;
   wire n_132_477;
   wire n_132_476;
   wire n_132_475;
   wire n_132_474;
   wire n_132_473;
   wire n_132_472;
   wire n_132_471;
   wire n_132_470;
   wire n_132_469;
   wire n_132_468;
   wire n_132_467;
   wire n_132_466;
   wire n_132_465;
   wire n_132_464;
   wire n_132_463;
   wire n_132_462;
   wire n_132_461;
   wire n_132_460;
   wire n_132_459;
   wire n_132_458;
   wire n_132_457;
   wire n_132_456;
   wire n_132_455;
   wire n_132_454;
   wire n_132_453;
   wire n_132_452;
   wire n_132_451;
   wire n_132_450;
   wire n_132_449;
   wire n_132_448;
   wire n_132_447;
   wire n_132_446;
   wire n_132_445;
   wire n_132_444;
   wire n_132_443;
   wire n_132_442;
   wire n_132_441;
   wire n_132_440;
   wire n_132_439;
   wire n_132_438;
   wire n_132_437;
   wire n_132_436;
   wire n_132_435;
   wire n_132_434;
   wire n_132_433;
   wire n_132_432;
   wire n_132_431;
   wire n_132_430;
   wire n_132_429;
   wire n_132_428;
   wire n_132_427;
   wire n_132_426;
   wire n_132_425;
   wire n_132_424;
   wire n_132_423;
   wire n_132_422;
   wire n_132_421;
   wire n_132_420;
   wire n_132_419;
   wire n_132_418;
   wire n_132_417;
   wire n_132_416;
   wire n_132_415;
   wire n_132_414;
   wire n_132_413;
   wire n_132_412;
   wire n_132_411;
   wire n_132_410;
   wire n_132_409;
   wire n_132_408;
   wire n_132_407;
   wire n_132_406;
   wire n_132_405;
   wire n_132_404;
   wire n_132_403;
   wire n_132_402;
   wire n_132_401;
   wire n_132_400;
   wire n_132_399;
   wire n_132_398;
   wire n_132_397;
   wire n_132_396;
   wire n_132_395;
   wire n_132_394;
   wire n_132_393;
   wire n_132_392;
   wire n_132_391;
   wire n_132_390;
   wire n_132_389;
   wire n_132_388;
   wire n_132_387;
   wire n_132_386;
   wire n_132_385;
   wire n_132_384;
   wire n_132_383;
   wire n_132_382;
   wire n_132_381;
   wire n_132_380;
   wire n_132_379;
   wire n_132_378;
   wire n_132_377;
   wire n_132_376;
   wire n_132_375;
   wire n_132_374;
   wire n_132_373;
   wire n_132_372;
   wire n_132_371;
   wire n_132_370;
   wire n_132_369;
   wire n_132_368;
   wire n_132_367;
   wire n_132_366;
   wire n_132_365;
   wire n_132_364;
   wire n_132_363;
   wire n_132_362;
   wire n_132_361;
   wire n_132_360;
   wire n_132_359;
   wire n_132_358;
   wire n_132_357;
   wire n_132_356;
   wire n_132_355;
   wire n_132_354;
   wire n_132_353;
   wire n_132_352;
   wire n_132_351;
   wire n_132_350;
   wire n_132_349;
   wire n_132_348;
   wire n_132_347;
   wire n_132_346;
   wire n_132_345;
   wire n_132_344;
   wire n_132_343;
   wire n_132_342;
   wire n_132_341;
   wire n_132_340;
   wire n_132_339;
   wire n_132_338;
   wire n_132_337;
   wire n_132_336;
   wire n_132_335;
   wire n_132_334;
   wire n_132_333;
   wire n_132_332;
   wire n_132_331;
   wire n_132_330;
   wire n_132_329;
   wire n_132_328;
   wire n_132_327;
   wire n_132_326;
   wire n_132_325;
   wire n_132_324;
   wire n_132_323;
   wire n_132_322;
   wire n_132_321;
   wire n_132_320;
   wire n_132_319;
   wire n_132_318;
   wire n_132_317;
   wire n_132_316;
   wire n_132_315;
   wire n_132_314;
   wire n_132_313;
   wire n_132_312;
   wire n_132_311;
   wire n_132_310;
   wire n_132_309;
   wire n_132_308;
   wire n_132_307;
   wire n_132_306;
   wire n_132_305;
   wire n_132_304;
   wire n_132_303;
   wire n_132_302;
   wire n_132_301;
   wire n_132_300;
   wire n_132_299;
   wire n_132_298;
   wire n_132_297;
   wire n_132_296;
   wire n_132_295;
   wire n_132_294;
   wire n_132_293;
   wire n_132_292;
   wire n_132_291;
   wire n_132_290;
   wire n_132_289;
   wire n_132_288;
   wire n_132_287;
   wire n_132_286;
   wire n_132_285;
   wire n_132_284;
   wire n_132_283;
   wire n_132_282;
   wire n_132_281;
   wire n_132_280;
   wire n_132_279;
   wire n_132_278;
   wire n_132_277;
   wire n_132_276;
   wire n_132_275;
   wire n_132_274;
   wire n_132_273;
   wire n_132_272;
   wire n_132_271;
   wire n_132_270;
   wire n_132_269;
   wire n_132_268;
   wire n_132_267;
   wire n_132_266;
   wire n_132_265;
   wire n_132_264;
   wire n_132_263;
   wire n_132_262;
   wire n_132_261;
   wire n_132_260;
   wire n_132_259;
   wire n_132_258;
   wire n_132_257;
   wire n_132_256;
   wire n_132_255;
   wire n_132_254;
   wire n_132_253;
   wire n_132_252;
   wire n_132_251;
   wire n_132_250;
   wire n_132_249;
   wire n_132_248;
   wire n_132_247;
   wire n_132_246;
   wire n_132_245;
   wire n_132_244;
   wire n_132_243;
   wire n_132_242;
   wire n_132_241;
   wire n_132_240;
   wire n_132_239;
   wire n_132_238;
   wire n_132_237;
   wire n_132_236;
   wire n_132_235;
   wire n_132_234;
   wire n_132_233;
   wire n_132_232;
   wire n_132_231;
   wire n_132_230;
   wire n_132_229;
   wire n_132_228;
   wire n_132_227;
   wire n_132_226;
   wire n_132_225;
   wire n_132_224;
   wire n_132_223;
   wire n_132_222;
   wire n_132_221;
   wire n_132_220;
   wire n_132_219;
   wire n_132_218;
   wire n_132_217;
   wire n_132_216;
   wire n_132_215;
   wire n_132_214;
   wire n_132_213;
   wire n_132_212;
   wire n_132_211;
   wire n_132_210;
   wire n_132_209;
   wire n_132_208;
   wire n_132_207;
   wire n_132_206;
   wire n_132_205;
   wire n_132_204;
   wire n_132_203;
   wire n_132_202;
   wire n_132_201;
   wire n_132_200;
   wire n_132_199;
   wire n_132_198;
   wire n_132_197;
   wire n_132_196;
   wire n_132_195;
   wire n_132_194;
   wire n_132_193;
   wire n_132_192;
   wire n_132_191;
   wire n_132_190;
   wire n_132_189;
   wire n_132_188;
   wire n_132_187;
   wire n_132_186;
   wire n_132_185;
   wire n_132_184;
   wire n_132_183;
   wire n_132_182;
   wire n_132_181;
   wire n_132_180;
   wire n_132_179;
   wire n_132_178;
   wire n_132_177;
   wire n_132_176;
   wire n_132_175;
   wire n_132_174;
   wire n_132_173;
   wire n_132_172;
   wire n_132_171;
   wire n_132_170;
   wire n_132_169;
   wire n_132_168;
   wire n_132_167;
   wire n_132_166;
   wire n_132_165;
   wire n_132_164;
   wire n_132_163;
   wire n_132_162;
   wire n_132_161;
   wire n_132_160;
   wire n_132_159;
   wire n_132_158;
   wire n_132_157;
   wire n_132_156;
   wire n_132_155;
   wire n_132_154;
   wire n_132_153;
   wire n_132_152;
   wire n_132_151;
   wire n_132_150;
   wire n_132_149;
   wire n_132_148;
   wire n_132_147;
   wire n_132_146;
   wire n_132_145;
   wire n_132_144;
   wire n_132_143;
   wire n_132_142;
   wire n_132_141;
   wire n_132_140;
   wire n_132_139;
   wire n_132_138;
   wire n_132_137;
   wire n_132_136;
   wire n_132_135;
   wire n_132_134;
   wire n_132_133;
   wire n_132_132;
   wire n_132_131;
   wire n_132_130;
   wire n_132_129;
   wire n_132_128;
   wire n_132_127;
   wire n_132_126;
   wire n_132_125;
   wire n_132_124;
   wire n_132_123;
   wire n_132_122;
   wire n_132_121;
   wire n_132_120;
   wire n_132_119;
   wire n_132_118;
   wire n_132_117;
   wire n_132_116;
   wire n_132_115;
   wire n_132_114;
   wire n_132_113;
   wire n_132_112;
   wire n_132_111;
   wire n_132_110;
   wire n_132_109;
   wire n_132_108;
   wire n_132_107;
   wire n_132_106;
   wire n_132_105;
   wire n_132_104;
   wire n_132_103;
   wire n_132_102;
   wire n_132_101;
   wire n_132_100;
   wire n_132_99;
   wire n_132_98;
   wire n_132_97;
   wire n_132_96;
   wire n_132_95;
   wire n_132_94;
   wire n_132_93;
   wire n_132_92;
   wire n_132_91;
   wire n_132_90;
   wire n_132_89;
   wire n_132_88;
   wire n_132_87;
   wire n_132_86;
   wire n_132_85;
   wire n_132_84;
   wire n_132_83;
   wire n_132_82;
   wire n_132_81;
   wire n_132_80;
   wire n_132_79;
   wire n_132_78;
   wire n_132_77;
   wire n_132_76;
   wire n_132_75;
   wire n_132_74;
   wire n_132_73;
   wire n_132_72;
   wire n_132_71;
   wire n_132_70;
   wire n_132_69;
   wire n_132_68;
   wire n_132_67;
   wire n_132_66;
   wire n_132_65;
   wire n_132_64;
   wire n_132_63;
   wire n_132_62;
   wire n_132_61;
   wire n_132_60;
   wire n_132_59;
   wire n_132_58;
   wire n_132_57;
   wire n_132_56;
   wire n_132_55;
   wire n_132_54;
   wire n_132_53;
   wire n_132_52;
   wire n_132_51;
   wire n_132_50;
   wire n_132_49;
   wire n_132_48;
   wire n_132_47;
   wire n_132_46;
   wire n_132_45;
   wire n_132_44;
   wire n_132_43;
   wire n_132_42;
   wire n_132_41;
   wire n_132_40;
   wire n_132_39;
   wire n_132_38;
   wire n_132_37;
   wire n_132_36;
   wire n_132_35;
   wire n_132_34;
   wire n_132_33;
   wire n_132_32;
   wire n_132_31;
   wire n_132_30;
   wire n_132_29;
   wire n_132_28;
   wire n_132_27;
   wire n_132_26;
   wire n_132_25;
   wire n_132_24;
   wire n_132_23;
   wire n_132_22;
   wire n_132_21;
   wire n_132_20;
   wire n_132_19;
   wire n_132_18;
   wire n_132_17;
   wire n_132_16;
   wire n_132_15;
   wire n_132_14;
   wire n_132_13;
   wire n_132_12;
   wire n_132_11;
   wire n_132_10;
   wire n_132_9;
   wire n_132_8;
   wire n_132_7;
   wire n_132_6;
   wire n_132_5;
   wire n_132_4;
   wire n_132_3;
   wire n_132_2;
   wire n_132_1;
   wire n_132_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0;
   wire n_0_0_38;
   wire n_0_1;
   wire n_0_0_39;
   wire n_0_62;
   wire n_0_0_40;
   wire n_0_61;
   wire n_0_0_41;
   wire n_0_60;
   wire n_0_0_42;
   wire n_0_59;
   wire n_0_0_43;
   wire n_0_58;
   wire n_0_0_44;
   wire n_0_57;
   wire n_0_0_45;
   wire n_0_56;
   wire n_0_0_46;
   wire n_0_55;
   wire n_0_0_47;
   wire n_0_54;
   wire n_0_0_48;
   wire n_0_53;
   wire n_0_0_49;
   wire n_0_52;
   wire n_0_0_50;
   wire n_0_51;
   wire n_0_0_51;
   wire n_0_50;
   wire n_0_0_52;
   wire n_0_49;
   wire n_0_0_53;
   wire n_0_48;
   wire n_0_0_54;
   wire n_0_47;
   wire n_0_0_55;
   wire n_0_46;
   wire n_0_0_56;
   wire n_0_45;
   wire n_0_0_57;
   wire n_0_44;
   wire n_0_0_58;
   wire n_0_43;
   wire n_0_0_59;
   wire n_0_42;
   wire n_0_0_60;
   wire n_0_41;
   wire n_0_0_61;
   wire n_0_40;
   wire n_0_0_62;
   wire n_0_39;
   wire n_0_0_63;
   wire n_0_38;
   wire n_0_0_64;
   wire n_0_37;
   wire n_0_0_65;
   wire n_0_36;
   wire n_0_0_66;
   wire n_0_35;
   wire n_0_0_67;
   wire n_0_34;
   wire n_0_0_68;
   wire n_0_33;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire read;
   wire n_1_3;
   wire [9:0]count;
   wire n_1_0;
   wire n_1_1;
   wire n_1_0_0;
   wire n_1_0_1;
   wire n_1_0_2;
   wire n_1_0_3;
   wire n_1_2;
   wire n_1_0_4;

   assign o_ready = 1'b1;

   DFF_X1 \o_buffer_reg[118][15]  (.D(n_123_959), .CK(n_120), .Q(
      \o_buffer[118] [15]), .QN());
   DFF_X1 \o_buffer_reg[118][14]  (.D(n_123_958), .CK(n_120), .Q(
      \o_buffer[118] [14]), .QN());
   DFF_X1 \o_buffer_reg[118][13]  (.D(n_123_957), .CK(n_120), .Q(
      \o_buffer[118] [13]), .QN());
   DFF_X1 \o_buffer_reg[118][12]  (.D(n_123_956), .CK(n_120), .Q(
      \o_buffer[118] [12]), .QN());
   DFF_X1 \o_buffer_reg[118][11]  (.D(n_123_955), .CK(n_120), .Q(
      \o_buffer[118] [11]), .QN());
   DFF_X1 \o_buffer_reg[118][10]  (.D(n_123_954), .CK(n_120), .Q(
      \o_buffer[118] [10]), .QN());
   DFF_X1 \o_buffer_reg[118][9]  (.D(n_123_953), .CK(n_120), .Q(
      \o_buffer[118] [9]), .QN());
   DFF_X1 \o_buffer_reg[118][8]  (.D(n_123_952), .CK(n_120), .Q(
      \o_buffer[118] [8]), .QN());
   DFF_X1 \o_buffer_reg[118][7]  (.D(n_123_951), .CK(n_120), .Q(
      \o_buffer[118] [7]), .QN());
   DFF_X1 \o_buffer_reg[118][6]  (.D(n_123_950), .CK(n_120), .Q(
      \o_buffer[118] [6]), .QN());
   DFF_X1 \o_buffer_reg[118][5]  (.D(n_123_949), .CK(n_120), .Q(
      \o_buffer[118] [5]), .QN());
   DFF_X1 \o_buffer_reg[118][4]  (.D(n_123_948), .CK(n_120), .Q(
      \o_buffer[118] [4]), .QN());
   DFF_X1 \o_buffer_reg[118][3]  (.D(n_123_947), .CK(n_120), .Q(
      \o_buffer[118] [3]), .QN());
   DFF_X1 \o_buffer_reg[118][2]  (.D(n_123_946), .CK(n_120), .Q(
      \o_buffer[118] [2]), .QN());
   DFF_X1 \o_buffer_reg[118][1]  (.D(n_123_945), .CK(n_120), .Q(
      \o_buffer[118] [1]), .QN());
   DFF_X1 \o_buffer_reg[118][0]  (.D(n_123_944), .CK(n_120), .Q(
      \o_buffer[118] [0]), .QN());
   DFF_X1 \o_buffer_reg[117][15]  (.D(n_123_943), .CK(n_120), .Q(
      \o_buffer[117] [15]), .QN());
   DFF_X1 \o_buffer_reg[117][14]  (.D(n_123_942), .CK(n_120), .Q(
      \o_buffer[117] [14]), .QN());
   DFF_X1 \o_buffer_reg[117][13]  (.D(n_123_941), .CK(n_120), .Q(
      \o_buffer[117] [13]), .QN());
   DFF_X1 \o_buffer_reg[117][12]  (.D(n_123_940), .CK(n_120), .Q(
      \o_buffer[117] [12]), .QN());
   DFF_X1 \o_buffer_reg[117][11]  (.D(n_123_939), .CK(n_120), .Q(
      \o_buffer[117] [11]), .QN());
   DFF_X1 \o_buffer_reg[117][10]  (.D(n_123_938), .CK(n_120), .Q(
      \o_buffer[117] [10]), .QN());
   DFF_X1 \o_buffer_reg[117][9]  (.D(n_123_937), .CK(n_120), .Q(
      \o_buffer[117] [9]), .QN());
   DFF_X1 \o_buffer_reg[117][8]  (.D(n_123_936), .CK(n_120), .Q(
      \o_buffer[117] [8]), .QN());
   DFF_X1 \o_buffer_reg[117][7]  (.D(n_123_935), .CK(n_120), .Q(
      \o_buffer[117] [7]), .QN());
   DFF_X1 \o_buffer_reg[117][6]  (.D(n_123_934), .CK(n_120), .Q(
      \o_buffer[117] [6]), .QN());
   DFF_X1 \o_buffer_reg[117][5]  (.D(n_123_933), .CK(n_120), .Q(
      \o_buffer[117] [5]), .QN());
   DFF_X1 \o_buffer_reg[117][4]  (.D(n_123_932), .CK(n_120), .Q(
      \o_buffer[117] [4]), .QN());
   DFF_X1 \o_buffer_reg[117][3]  (.D(n_123_931), .CK(n_120), .Q(
      \o_buffer[117] [3]), .QN());
   DFF_X1 \o_buffer_reg[117][2]  (.D(n_123_930), .CK(n_120), .Q(
      \o_buffer[117] [2]), .QN());
   DFF_X1 \o_buffer_reg[117][1]  (.D(n_123_929), .CK(n_120), .Q(
      \o_buffer[117] [1]), .QN());
   DFF_X1 \o_buffer_reg[117][0]  (.D(n_123_928), .CK(n_120), .Q(
      \o_buffer[117] [0]), .QN());
   DFF_X1 \o_buffer_reg[116][15]  (.D(n_123_927), .CK(n_120), .Q(
      \o_buffer[116] [15]), .QN());
   DFF_X1 \o_buffer_reg[116][14]  (.D(n_123_926), .CK(n_120), .Q(
      \o_buffer[116] [14]), .QN());
   DFF_X1 \o_buffer_reg[116][13]  (.D(n_123_925), .CK(n_120), .Q(
      \o_buffer[116] [13]), .QN());
   DFF_X1 \o_buffer_reg[116][12]  (.D(n_123_924), .CK(n_120), .Q(
      \o_buffer[116] [12]), .QN());
   DFF_X1 \o_buffer_reg[116][11]  (.D(n_123_923), .CK(n_120), .Q(
      \o_buffer[116] [11]), .QN());
   DFF_X1 \o_buffer_reg[116][10]  (.D(n_123_922), .CK(n_120), .Q(
      \o_buffer[116] [10]), .QN());
   DFF_X1 \o_buffer_reg[116][9]  (.D(n_123_921), .CK(n_120), .Q(
      \o_buffer[116] [9]), .QN());
   DFF_X1 \o_buffer_reg[116][8]  (.D(n_123_920), .CK(n_120), .Q(
      \o_buffer[116] [8]), .QN());
   DFF_X1 \o_buffer_reg[116][7]  (.D(n_123_919), .CK(n_120), .Q(
      \o_buffer[116] [7]), .QN());
   DFF_X1 \o_buffer_reg[116][6]  (.D(n_123_918), .CK(n_120), .Q(
      \o_buffer[116] [6]), .QN());
   DFF_X1 \o_buffer_reg[116][5]  (.D(n_123_917), .CK(n_120), .Q(
      \o_buffer[116] [5]), .QN());
   DFF_X1 \o_buffer_reg[116][4]  (.D(n_123_916), .CK(n_120), .Q(
      \o_buffer[116] [4]), .QN());
   DFF_X1 \o_buffer_reg[116][3]  (.D(n_123_915), .CK(n_120), .Q(
      \o_buffer[116] [3]), .QN());
   DFF_X1 \o_buffer_reg[116][2]  (.D(n_123_914), .CK(n_120), .Q(
      \o_buffer[116] [2]), .QN());
   DFF_X1 \o_buffer_reg[116][1]  (.D(n_123_913), .CK(n_120), .Q(
      \o_buffer[116] [1]), .QN());
   DFF_X1 \o_buffer_reg[116][0]  (.D(n_123_912), .CK(n_120), .Q(
      \o_buffer[116] [0]), .QN());
   DFF_X1 \o_buffer_reg[115][15]  (.D(n_123_911), .CK(n_120), .Q(
      \o_buffer[115] [15]), .QN());
   DFF_X1 \o_buffer_reg[115][14]  (.D(n_123_910), .CK(n_120), .Q(
      \o_buffer[115] [14]), .QN());
   DFF_X1 \o_buffer_reg[115][13]  (.D(n_123_909), .CK(n_120), .Q(
      \o_buffer[115] [13]), .QN());
   DFF_X1 \o_buffer_reg[115][12]  (.D(n_123_908), .CK(n_120), .Q(
      \o_buffer[115] [12]), .QN());
   DFF_X1 \o_buffer_reg[115][11]  (.D(n_123_907), .CK(n_120), .Q(
      \o_buffer[115] [11]), .QN());
   DFF_X1 \o_buffer_reg[115][10]  (.D(n_123_906), .CK(n_120), .Q(
      \o_buffer[115] [10]), .QN());
   DFF_X1 \o_buffer_reg[115][9]  (.D(n_123_905), .CK(n_120), .Q(
      \o_buffer[115] [9]), .QN());
   DFF_X1 \o_buffer_reg[115][8]  (.D(n_123_904), .CK(n_120), .Q(
      \o_buffer[115] [8]), .QN());
   DFF_X1 \o_buffer_reg[115][7]  (.D(n_123_903), .CK(n_120), .Q(
      \o_buffer[115] [7]), .QN());
   DFF_X1 \o_buffer_reg[115][6]  (.D(n_123_902), .CK(n_120), .Q(
      \o_buffer[115] [6]), .QN());
   DFF_X1 \o_buffer_reg[115][5]  (.D(n_123_901), .CK(n_120), .Q(
      \o_buffer[115] [5]), .QN());
   DFF_X1 \o_buffer_reg[115][4]  (.D(n_123_900), .CK(n_120), .Q(
      \o_buffer[115] [4]), .QN());
   DFF_X1 \o_buffer_reg[115][3]  (.D(n_123_899), .CK(n_120), .Q(
      \o_buffer[115] [3]), .QN());
   DFF_X1 \o_buffer_reg[115][2]  (.D(n_123_898), .CK(n_120), .Q(
      \o_buffer[115] [2]), .QN());
   DFF_X1 \o_buffer_reg[115][1]  (.D(n_123_897), .CK(n_120), .Q(
      \o_buffer[115] [1]), .QN());
   DFF_X1 \o_buffer_reg[115][0]  (.D(n_123_896), .CK(n_120), .Q(
      \o_buffer[115] [0]), .QN());
   DFF_X1 \o_buffer_reg[114][15]  (.D(n_123_895), .CK(n_120), .Q(
      \o_buffer[114] [15]), .QN());
   DFF_X1 \o_buffer_reg[114][14]  (.D(n_123_894), .CK(n_120), .Q(
      \o_buffer[114] [14]), .QN());
   DFF_X1 \o_buffer_reg[114][13]  (.D(n_123_893), .CK(n_120), .Q(
      \o_buffer[114] [13]), .QN());
   DFF_X1 \o_buffer_reg[114][12]  (.D(n_123_892), .CK(n_120), .Q(
      \o_buffer[114] [12]), .QN());
   DFF_X1 \o_buffer_reg[114][11]  (.D(n_123_891), .CK(n_120), .Q(
      \o_buffer[114] [11]), .QN());
   DFF_X1 \o_buffer_reg[114][10]  (.D(n_123_890), .CK(n_120), .Q(
      \o_buffer[114] [10]), .QN());
   DFF_X1 \o_buffer_reg[114][9]  (.D(n_123_889), .CK(n_120), .Q(
      \o_buffer[114] [9]), .QN());
   DFF_X1 \o_buffer_reg[114][8]  (.D(n_123_888), .CK(n_120), .Q(
      \o_buffer[114] [8]), .QN());
   DFF_X1 \o_buffer_reg[114][7]  (.D(n_123_887), .CK(n_120), .Q(
      \o_buffer[114] [7]), .QN());
   DFF_X1 \o_buffer_reg[114][6]  (.D(n_123_886), .CK(n_120), .Q(
      \o_buffer[114] [6]), .QN());
   DFF_X1 \o_buffer_reg[114][5]  (.D(n_123_885), .CK(n_120), .Q(
      \o_buffer[114] [5]), .QN());
   DFF_X1 \o_buffer_reg[114][4]  (.D(n_123_884), .CK(n_120), .Q(
      \o_buffer[114] [4]), .QN());
   DFF_X1 \o_buffer_reg[114][3]  (.D(n_123_883), .CK(n_120), .Q(
      \o_buffer[114] [3]), .QN());
   DFF_X1 \o_buffer_reg[114][2]  (.D(n_123_882), .CK(n_120), .Q(
      \o_buffer[114] [2]), .QN());
   DFF_X1 \o_buffer_reg[114][1]  (.D(n_123_881), .CK(n_120), .Q(
      \o_buffer[114] [1]), .QN());
   DFF_X1 \o_buffer_reg[114][0]  (.D(n_123_880), .CK(n_120), .Q(
      \o_buffer[114] [0]), .QN());
   DFF_X1 \o_buffer_reg[113][15]  (.D(n_123_879), .CK(n_120), .Q(
      \o_buffer[113] [15]), .QN());
   DFF_X1 \o_buffer_reg[113][14]  (.D(n_123_878), .CK(n_120), .Q(
      \o_buffer[113] [14]), .QN());
   DFF_X1 \o_buffer_reg[113][13]  (.D(n_123_877), .CK(n_120), .Q(
      \o_buffer[113] [13]), .QN());
   DFF_X1 \o_buffer_reg[113][12]  (.D(n_123_876), .CK(n_120), .Q(
      \o_buffer[113] [12]), .QN());
   DFF_X1 \o_buffer_reg[113][11]  (.D(n_123_875), .CK(n_120), .Q(
      \o_buffer[113] [11]), .QN());
   DFF_X1 \o_buffer_reg[113][10]  (.D(n_123_874), .CK(n_120), .Q(
      \o_buffer[113] [10]), .QN());
   DFF_X1 \o_buffer_reg[113][9]  (.D(n_123_873), .CK(n_120), .Q(
      \o_buffer[113] [9]), .QN());
   DFF_X1 \o_buffer_reg[113][8]  (.D(n_123_872), .CK(n_120), .Q(
      \o_buffer[113] [8]), .QN());
   DFF_X1 \o_buffer_reg[113][7]  (.D(n_123_871), .CK(n_120), .Q(
      \o_buffer[113] [7]), .QN());
   DFF_X1 \o_buffer_reg[113][6]  (.D(n_123_870), .CK(n_120), .Q(
      \o_buffer[113] [6]), .QN());
   DFF_X1 \o_buffer_reg[113][5]  (.D(n_123_869), .CK(n_120), .Q(
      \o_buffer[113] [5]), .QN());
   DFF_X1 \o_buffer_reg[113][4]  (.D(n_123_868), .CK(n_120), .Q(
      \o_buffer[113] [4]), .QN());
   DFF_X1 \o_buffer_reg[113][3]  (.D(n_123_867), .CK(n_120), .Q(
      \o_buffer[113] [3]), .QN());
   DFF_X1 \o_buffer_reg[113][2]  (.D(n_123_866), .CK(n_120), .Q(
      \o_buffer[113] [2]), .QN());
   DFF_X1 \o_buffer_reg[113][1]  (.D(n_123_865), .CK(n_120), .Q(
      \o_buffer[113] [1]), .QN());
   DFF_X1 \o_buffer_reg[113][0]  (.D(n_123_864), .CK(n_120), .Q(
      \o_buffer[113] [0]), .QN());
   DFF_X1 \o_buffer_reg[112][15]  (.D(n_123_863), .CK(n_120), .Q(
      \o_buffer[112] [15]), .QN());
   DFF_X1 \o_buffer_reg[112][14]  (.D(n_123_862), .CK(n_120), .Q(
      \o_buffer[112] [14]), .QN());
   DFF_X1 \o_buffer_reg[112][13]  (.D(n_123_861), .CK(n_120), .Q(
      \o_buffer[112] [13]), .QN());
   DFF_X1 \o_buffer_reg[112][12]  (.D(n_123_860), .CK(n_120), .Q(
      \o_buffer[112] [12]), .QN());
   DFF_X1 \o_buffer_reg[112][11]  (.D(n_123_859), .CK(n_120), .Q(
      \o_buffer[112] [11]), .QN());
   DFF_X1 \o_buffer_reg[112][10]  (.D(n_123_858), .CK(n_120), .Q(
      \o_buffer[112] [10]), .QN());
   DFF_X1 \o_buffer_reg[112][9]  (.D(n_123_857), .CK(n_120), .Q(
      \o_buffer[112] [9]), .QN());
   DFF_X1 \o_buffer_reg[112][8]  (.D(n_123_856), .CK(n_120), .Q(
      \o_buffer[112] [8]), .QN());
   DFF_X1 \o_buffer_reg[112][7]  (.D(n_123_855), .CK(n_120), .Q(
      \o_buffer[112] [7]), .QN());
   DFF_X1 \o_buffer_reg[112][6]  (.D(n_123_854), .CK(n_120), .Q(
      \o_buffer[112] [6]), .QN());
   DFF_X1 \o_buffer_reg[112][5]  (.D(n_123_853), .CK(n_120), .Q(
      \o_buffer[112] [5]), .QN());
   DFF_X1 \o_buffer_reg[112][4]  (.D(n_123_852), .CK(n_120), .Q(
      \o_buffer[112] [4]), .QN());
   DFF_X1 \o_buffer_reg[112][3]  (.D(n_123_851), .CK(n_120), .Q(
      \o_buffer[112] [3]), .QN());
   DFF_X1 \o_buffer_reg[112][2]  (.D(n_123_850), .CK(n_120), .Q(
      \o_buffer[112] [2]), .QN());
   DFF_X1 \o_buffer_reg[112][1]  (.D(n_123_849), .CK(n_120), .Q(
      \o_buffer[112] [1]), .QN());
   DFF_X1 \o_buffer_reg[112][0]  (.D(n_123_848), .CK(n_120), .Q(
      \o_buffer[112] [0]), .QN());
   DFF_X1 \o_buffer_reg[111][15]  (.D(n_123_847), .CK(n_120), .Q(
      \o_buffer[111] [15]), .QN());
   DFF_X1 \o_buffer_reg[111][14]  (.D(n_123_846), .CK(n_120), .Q(
      \o_buffer[111] [14]), .QN());
   DFF_X1 \o_buffer_reg[111][13]  (.D(n_123_845), .CK(n_120), .Q(
      \o_buffer[111] [13]), .QN());
   DFF_X1 \o_buffer_reg[111][12]  (.D(n_123_844), .CK(n_120), .Q(
      \o_buffer[111] [12]), .QN());
   DFF_X1 \o_buffer_reg[111][11]  (.D(n_123_843), .CK(n_120), .Q(
      \o_buffer[111] [11]), .QN());
   DFF_X1 \o_buffer_reg[111][10]  (.D(n_123_842), .CK(n_120), .Q(
      \o_buffer[111] [10]), .QN());
   DFF_X1 \o_buffer_reg[111][9]  (.D(n_123_841), .CK(n_120), .Q(
      \o_buffer[111] [9]), .QN());
   DFF_X1 \o_buffer_reg[111][8]  (.D(n_123_840), .CK(n_120), .Q(
      \o_buffer[111] [8]), .QN());
   DFF_X1 \o_buffer_reg[111][7]  (.D(n_123_839), .CK(n_120), .Q(
      \o_buffer[111] [7]), .QN());
   DFF_X1 \o_buffer_reg[111][6]  (.D(n_123_838), .CK(n_120), .Q(
      \o_buffer[111] [6]), .QN());
   DFF_X1 \o_buffer_reg[111][5]  (.D(n_123_837), .CK(n_120), .Q(
      \o_buffer[111] [5]), .QN());
   DFF_X1 \o_buffer_reg[111][4]  (.D(n_123_836), .CK(n_120), .Q(
      \o_buffer[111] [4]), .QN());
   DFF_X1 \o_buffer_reg[111][3]  (.D(n_123_835), .CK(n_120), .Q(
      \o_buffer[111] [3]), .QN());
   DFF_X1 \o_buffer_reg[111][2]  (.D(n_123_834), .CK(n_120), .Q(
      \o_buffer[111] [2]), .QN());
   DFF_X1 \o_buffer_reg[111][1]  (.D(n_123_833), .CK(n_120), .Q(
      \o_buffer[111] [1]), .QN());
   DFF_X1 \o_buffer_reg[111][0]  (.D(n_123_832), .CK(n_120), .Q(
      \o_buffer[111] [0]), .QN());
   DFF_X1 \o_buffer_reg[110][15]  (.D(n_123_831), .CK(n_120), .Q(
      \o_buffer[110] [15]), .QN());
   DFF_X1 \o_buffer_reg[110][14]  (.D(n_123_830), .CK(n_120), .Q(
      \o_buffer[110] [14]), .QN());
   DFF_X1 \o_buffer_reg[110][13]  (.D(n_123_829), .CK(n_120), .Q(
      \o_buffer[110] [13]), .QN());
   DFF_X1 \o_buffer_reg[110][12]  (.D(n_123_828), .CK(n_120), .Q(
      \o_buffer[110] [12]), .QN());
   DFF_X1 \o_buffer_reg[110][11]  (.D(n_123_827), .CK(n_120), .Q(
      \o_buffer[110] [11]), .QN());
   DFF_X1 \o_buffer_reg[110][10]  (.D(n_123_826), .CK(n_120), .Q(
      \o_buffer[110] [10]), .QN());
   DFF_X1 \o_buffer_reg[110][9]  (.D(n_123_825), .CK(n_120), .Q(
      \o_buffer[110] [9]), .QN());
   DFF_X1 \o_buffer_reg[110][8]  (.D(n_123_824), .CK(n_120), .Q(
      \o_buffer[110] [8]), .QN());
   DFF_X1 \o_buffer_reg[110][7]  (.D(n_123_823), .CK(n_120), .Q(
      \o_buffer[110] [7]), .QN());
   DFF_X1 \o_buffer_reg[110][6]  (.D(n_123_822), .CK(n_120), .Q(
      \o_buffer[110] [6]), .QN());
   DFF_X1 \o_buffer_reg[110][5]  (.D(n_123_821), .CK(n_120), .Q(
      \o_buffer[110] [5]), .QN());
   DFF_X1 \o_buffer_reg[110][4]  (.D(n_123_820), .CK(n_120), .Q(
      \o_buffer[110] [4]), .QN());
   DFF_X1 \o_buffer_reg[110][3]  (.D(n_123_819), .CK(n_120), .Q(
      \o_buffer[110] [3]), .QN());
   DFF_X1 \o_buffer_reg[110][2]  (.D(n_123_818), .CK(n_120), .Q(
      \o_buffer[110] [2]), .QN());
   DFF_X1 \o_buffer_reg[110][1]  (.D(n_123_817), .CK(n_120), .Q(
      \o_buffer[110] [1]), .QN());
   DFF_X1 \o_buffer_reg[110][0]  (.D(n_123_816), .CK(n_120), .Q(
      \o_buffer[110] [0]), .QN());
   DFF_X1 \o_buffer_reg[109][15]  (.D(n_123_815), .CK(n_120), .Q(
      \o_buffer[109] [15]), .QN());
   DFF_X1 \o_buffer_reg[109][14]  (.D(n_123_814), .CK(n_120), .Q(
      \o_buffer[109] [14]), .QN());
   DFF_X1 \o_buffer_reg[109][13]  (.D(n_123_813), .CK(n_120), .Q(
      \o_buffer[109] [13]), .QN());
   DFF_X1 \o_buffer_reg[109][12]  (.D(n_123_812), .CK(n_120), .Q(
      \o_buffer[109] [12]), .QN());
   DFF_X1 \o_buffer_reg[109][11]  (.D(n_123_811), .CK(n_120), .Q(
      \o_buffer[109] [11]), .QN());
   DFF_X1 \o_buffer_reg[109][10]  (.D(n_123_810), .CK(n_120), .Q(
      \o_buffer[109] [10]), .QN());
   DFF_X1 \o_buffer_reg[109][9]  (.D(n_123_809), .CK(n_120), .Q(
      \o_buffer[109] [9]), .QN());
   DFF_X1 \o_buffer_reg[109][8]  (.D(n_123_808), .CK(n_120), .Q(
      \o_buffer[109] [8]), .QN());
   DFF_X1 \o_buffer_reg[109][7]  (.D(n_123_807), .CK(n_120), .Q(
      \o_buffer[109] [7]), .QN());
   DFF_X1 \o_buffer_reg[109][6]  (.D(n_123_806), .CK(n_120), .Q(
      \o_buffer[109] [6]), .QN());
   DFF_X1 \o_buffer_reg[109][5]  (.D(n_123_805), .CK(n_120), .Q(
      \o_buffer[109] [5]), .QN());
   DFF_X1 \o_buffer_reg[109][4]  (.D(n_123_804), .CK(n_120), .Q(
      \o_buffer[109] [4]), .QN());
   DFF_X1 \o_buffer_reg[109][3]  (.D(n_123_803), .CK(n_120), .Q(
      \o_buffer[109] [3]), .QN());
   DFF_X1 \o_buffer_reg[109][2]  (.D(n_123_802), .CK(n_120), .Q(
      \o_buffer[109] [2]), .QN());
   DFF_X1 \o_buffer_reg[109][1]  (.D(n_123_801), .CK(n_120), .Q(
      \o_buffer[109] [1]), .QN());
   DFF_X1 \o_buffer_reg[109][0]  (.D(n_123_800), .CK(n_120), .Q(
      \o_buffer[109] [0]), .QN());
   DFF_X1 \o_buffer_reg[108][15]  (.D(n_123_799), .CK(n_120), .Q(
      \o_buffer[108] [15]), .QN());
   DFF_X1 \o_buffer_reg[108][14]  (.D(n_123_798), .CK(n_120), .Q(
      \o_buffer[108] [14]), .QN());
   DFF_X1 \o_buffer_reg[108][13]  (.D(n_123_797), .CK(n_120), .Q(
      \o_buffer[108] [13]), .QN());
   DFF_X1 \o_buffer_reg[108][12]  (.D(n_123_796), .CK(n_120), .Q(
      \o_buffer[108] [12]), .QN());
   DFF_X1 \o_buffer_reg[108][11]  (.D(n_123_795), .CK(n_120), .Q(
      \o_buffer[108] [11]), .QN());
   DFF_X1 \o_buffer_reg[108][10]  (.D(n_123_794), .CK(n_120), .Q(
      \o_buffer[108] [10]), .QN());
   DFF_X1 \o_buffer_reg[108][9]  (.D(n_123_793), .CK(n_120), .Q(
      \o_buffer[108] [9]), .QN());
   DFF_X1 \o_buffer_reg[108][8]  (.D(n_123_792), .CK(n_120), .Q(
      \o_buffer[108] [8]), .QN());
   DFF_X1 \o_buffer_reg[108][7]  (.D(n_123_791), .CK(n_120), .Q(
      \o_buffer[108] [7]), .QN());
   DFF_X1 \o_buffer_reg[108][6]  (.D(n_123_790), .CK(n_120), .Q(
      \o_buffer[108] [6]), .QN());
   DFF_X1 \o_buffer_reg[108][5]  (.D(n_123_789), .CK(n_120), .Q(
      \o_buffer[108] [5]), .QN());
   DFF_X1 \o_buffer_reg[108][4]  (.D(n_123_788), .CK(n_120), .Q(
      \o_buffer[108] [4]), .QN());
   DFF_X1 \o_buffer_reg[108][3]  (.D(n_123_787), .CK(n_120), .Q(
      \o_buffer[108] [3]), .QN());
   DFF_X1 \o_buffer_reg[108][2]  (.D(n_123_786), .CK(n_120), .Q(
      \o_buffer[108] [2]), .QN());
   DFF_X1 \o_buffer_reg[108][1]  (.D(n_123_785), .CK(n_120), .Q(
      \o_buffer[108] [1]), .QN());
   DFF_X1 \o_buffer_reg[108][0]  (.D(n_123_784), .CK(n_120), .Q(
      \o_buffer[108] [0]), .QN());
   DFF_X1 \o_buffer_reg[107][15]  (.D(n_123_783), .CK(n_120), .Q(
      \o_buffer[107] [15]), .QN());
   DFF_X1 \o_buffer_reg[107][14]  (.D(n_123_782), .CK(n_120), .Q(
      \o_buffer[107] [14]), .QN());
   DFF_X1 \o_buffer_reg[107][13]  (.D(n_123_781), .CK(n_120), .Q(
      \o_buffer[107] [13]), .QN());
   DFF_X1 \o_buffer_reg[107][12]  (.D(n_123_780), .CK(n_120), .Q(
      \o_buffer[107] [12]), .QN());
   DFF_X1 \o_buffer_reg[107][11]  (.D(n_123_779), .CK(n_120), .Q(
      \o_buffer[107] [11]), .QN());
   DFF_X1 \o_buffer_reg[107][10]  (.D(n_123_778), .CK(n_120), .Q(
      \o_buffer[107] [10]), .QN());
   DFF_X1 \o_buffer_reg[107][9]  (.D(n_123_777), .CK(n_120), .Q(
      \o_buffer[107] [9]), .QN());
   DFF_X1 \o_buffer_reg[107][8]  (.D(n_123_776), .CK(n_120), .Q(
      \o_buffer[107] [8]), .QN());
   DFF_X1 \o_buffer_reg[107][7]  (.D(n_123_775), .CK(n_120), .Q(
      \o_buffer[107] [7]), .QN());
   DFF_X1 \o_buffer_reg[107][6]  (.D(n_123_774), .CK(n_120), .Q(
      \o_buffer[107] [6]), .QN());
   DFF_X1 \o_buffer_reg[107][5]  (.D(n_123_773), .CK(n_120), .Q(
      \o_buffer[107] [5]), .QN());
   DFF_X1 \o_buffer_reg[107][4]  (.D(n_123_772), .CK(n_120), .Q(
      \o_buffer[107] [4]), .QN());
   DFF_X1 \o_buffer_reg[107][3]  (.D(n_123_771), .CK(n_120), .Q(
      \o_buffer[107] [3]), .QN());
   DFF_X1 \o_buffer_reg[107][2]  (.D(n_123_770), .CK(n_120), .Q(
      \o_buffer[107] [2]), .QN());
   DFF_X1 \o_buffer_reg[107][1]  (.D(n_123_769), .CK(n_120), .Q(
      \o_buffer[107] [1]), .QN());
   DFF_X1 \o_buffer_reg[107][0]  (.D(n_123_768), .CK(n_120), .Q(
      \o_buffer[107] [0]), .QN());
   DFF_X1 \o_buffer_reg[106][15]  (.D(n_123_767), .CK(n_120), .Q(
      \o_buffer[106] [15]), .QN());
   DFF_X1 \o_buffer_reg[106][14]  (.D(n_123_766), .CK(n_120), .Q(
      \o_buffer[106] [14]), .QN());
   DFF_X1 \o_buffer_reg[106][13]  (.D(n_123_765), .CK(n_120), .Q(
      \o_buffer[106] [13]), .QN());
   DFF_X1 \o_buffer_reg[106][12]  (.D(n_123_764), .CK(n_120), .Q(
      \o_buffer[106] [12]), .QN());
   DFF_X1 \o_buffer_reg[106][11]  (.D(n_123_763), .CK(n_120), .Q(
      \o_buffer[106] [11]), .QN());
   DFF_X1 \o_buffer_reg[106][10]  (.D(n_123_762), .CK(n_120), .Q(
      \o_buffer[106] [10]), .QN());
   DFF_X1 \o_buffer_reg[106][9]  (.D(n_123_761), .CK(n_120), .Q(
      \o_buffer[106] [9]), .QN());
   DFF_X1 \o_buffer_reg[106][8]  (.D(n_123_760), .CK(n_120), .Q(
      \o_buffer[106] [8]), .QN());
   DFF_X1 \o_buffer_reg[106][7]  (.D(n_123_759), .CK(n_120), .Q(
      \o_buffer[106] [7]), .QN());
   DFF_X1 \o_buffer_reg[106][6]  (.D(n_123_758), .CK(n_120), .Q(
      \o_buffer[106] [6]), .QN());
   DFF_X1 \o_buffer_reg[106][5]  (.D(n_123_757), .CK(n_120), .Q(
      \o_buffer[106] [5]), .QN());
   DFF_X1 \o_buffer_reg[106][4]  (.D(n_123_756), .CK(n_120), .Q(
      \o_buffer[106] [4]), .QN());
   DFF_X1 \o_buffer_reg[106][3]  (.D(n_123_755), .CK(n_120), .Q(
      \o_buffer[106] [3]), .QN());
   DFF_X1 \o_buffer_reg[106][2]  (.D(n_123_754), .CK(n_120), .Q(
      \o_buffer[106] [2]), .QN());
   DFF_X1 \o_buffer_reg[106][1]  (.D(n_123_753), .CK(n_120), .Q(
      \o_buffer[106] [1]), .QN());
   DFF_X1 \o_buffer_reg[106][0]  (.D(n_123_752), .CK(n_120), .Q(
      \o_buffer[106] [0]), .QN());
   DFF_X1 \o_buffer_reg[105][15]  (.D(n_123_751), .CK(n_120), .Q(
      \o_buffer[105] [15]), .QN());
   DFF_X1 \o_buffer_reg[105][14]  (.D(n_123_750), .CK(n_120), .Q(
      \o_buffer[105] [14]), .QN());
   DFF_X1 \o_buffer_reg[105][13]  (.D(n_123_749), .CK(n_120), .Q(
      \o_buffer[105] [13]), .QN());
   DFF_X1 \o_buffer_reg[105][12]  (.D(n_123_748), .CK(n_120), .Q(
      \o_buffer[105] [12]), .QN());
   DFF_X1 \o_buffer_reg[105][11]  (.D(n_123_747), .CK(n_120), .Q(
      \o_buffer[105] [11]), .QN());
   DFF_X1 \o_buffer_reg[105][10]  (.D(n_123_746), .CK(n_120), .Q(
      \o_buffer[105] [10]), .QN());
   DFF_X1 \o_buffer_reg[105][9]  (.D(n_123_745), .CK(n_120), .Q(
      \o_buffer[105] [9]), .QN());
   DFF_X1 \o_buffer_reg[105][8]  (.D(n_123_744), .CK(n_120), .Q(
      \o_buffer[105] [8]), .QN());
   DFF_X1 \o_buffer_reg[105][7]  (.D(n_123_743), .CK(n_120), .Q(
      \o_buffer[105] [7]), .QN());
   DFF_X1 \o_buffer_reg[105][6]  (.D(n_123_742), .CK(n_120), .Q(
      \o_buffer[105] [6]), .QN());
   DFF_X1 \o_buffer_reg[105][5]  (.D(n_123_741), .CK(n_120), .Q(
      \o_buffer[105] [5]), .QN());
   DFF_X1 \o_buffer_reg[105][4]  (.D(n_123_740), .CK(n_120), .Q(
      \o_buffer[105] [4]), .QN());
   DFF_X1 \o_buffer_reg[105][3]  (.D(n_123_739), .CK(n_120), .Q(
      \o_buffer[105] [3]), .QN());
   DFF_X1 \o_buffer_reg[105][2]  (.D(n_123_738), .CK(n_120), .Q(
      \o_buffer[105] [2]), .QN());
   DFF_X1 \o_buffer_reg[105][1]  (.D(n_123_737), .CK(n_120), .Q(
      \o_buffer[105] [1]), .QN());
   DFF_X1 \o_buffer_reg[105][0]  (.D(n_123_736), .CK(n_120), .Q(
      \o_buffer[105] [0]), .QN());
   DFF_X1 \o_buffer_reg[104][15]  (.D(n_123_735), .CK(n_120), .Q(
      \o_buffer[104] [15]), .QN());
   DFF_X1 \o_buffer_reg[104][14]  (.D(n_123_734), .CK(n_120), .Q(
      \o_buffer[104] [14]), .QN());
   DFF_X1 \o_buffer_reg[104][13]  (.D(n_123_733), .CK(n_120), .Q(
      \o_buffer[104] [13]), .QN());
   DFF_X1 \o_buffer_reg[104][12]  (.D(n_123_732), .CK(n_120), .Q(
      \o_buffer[104] [12]), .QN());
   DFF_X1 \o_buffer_reg[104][11]  (.D(n_123_731), .CK(n_120), .Q(
      \o_buffer[104] [11]), .QN());
   DFF_X1 \o_buffer_reg[104][10]  (.D(n_123_730), .CK(n_120), .Q(
      \o_buffer[104] [10]), .QN());
   DFF_X1 \o_buffer_reg[104][9]  (.D(n_123_729), .CK(n_120), .Q(
      \o_buffer[104] [9]), .QN());
   DFF_X1 \o_buffer_reg[104][8]  (.D(n_123_728), .CK(n_120), .Q(
      \o_buffer[104] [8]), .QN());
   DFF_X1 \o_buffer_reg[104][7]  (.D(n_123_727), .CK(n_120), .Q(
      \o_buffer[104] [7]), .QN());
   DFF_X1 \o_buffer_reg[104][6]  (.D(n_123_726), .CK(n_120), .Q(
      \o_buffer[104] [6]), .QN());
   DFF_X1 \o_buffer_reg[104][5]  (.D(n_123_725), .CK(n_120), .Q(
      \o_buffer[104] [5]), .QN());
   DFF_X1 \o_buffer_reg[104][4]  (.D(n_123_724), .CK(n_120), .Q(
      \o_buffer[104] [4]), .QN());
   DFF_X1 \o_buffer_reg[104][3]  (.D(n_123_723), .CK(n_120), .Q(
      \o_buffer[104] [3]), .QN());
   DFF_X1 \o_buffer_reg[104][2]  (.D(n_123_722), .CK(n_120), .Q(
      \o_buffer[104] [2]), .QN());
   DFF_X1 \o_buffer_reg[104][1]  (.D(n_123_721), .CK(n_120), .Q(
      \o_buffer[104] [1]), .QN());
   DFF_X1 \o_buffer_reg[104][0]  (.D(n_123_720), .CK(n_120), .Q(
      \o_buffer[104] [0]), .QN());
   DFF_X1 \o_buffer_reg[103][15]  (.D(n_123_719), .CK(n_120), .Q(
      \o_buffer[103] [15]), .QN());
   DFF_X1 \o_buffer_reg[103][14]  (.D(n_123_718), .CK(n_120), .Q(
      \o_buffer[103] [14]), .QN());
   DFF_X1 \o_buffer_reg[103][13]  (.D(n_123_717), .CK(n_120), .Q(
      \o_buffer[103] [13]), .QN());
   DFF_X1 \o_buffer_reg[103][12]  (.D(n_123_716), .CK(n_120), .Q(
      \o_buffer[103] [12]), .QN());
   DFF_X1 \o_buffer_reg[103][11]  (.D(n_123_715), .CK(n_120), .Q(
      \o_buffer[103] [11]), .QN());
   DFF_X1 \o_buffer_reg[103][10]  (.D(n_123_714), .CK(n_120), .Q(
      \o_buffer[103] [10]), .QN());
   DFF_X1 \o_buffer_reg[103][9]  (.D(n_123_713), .CK(n_120), .Q(
      \o_buffer[103] [9]), .QN());
   DFF_X1 \o_buffer_reg[103][8]  (.D(n_123_712), .CK(n_120), .Q(
      \o_buffer[103] [8]), .QN());
   DFF_X1 \o_buffer_reg[103][7]  (.D(n_123_711), .CK(n_120), .Q(
      \o_buffer[103] [7]), .QN());
   DFF_X1 \o_buffer_reg[103][6]  (.D(n_123_710), .CK(n_120), .Q(
      \o_buffer[103] [6]), .QN());
   DFF_X1 \o_buffer_reg[103][5]  (.D(n_123_709), .CK(n_120), .Q(
      \o_buffer[103] [5]), .QN());
   DFF_X1 \o_buffer_reg[103][4]  (.D(n_123_708), .CK(n_120), .Q(
      \o_buffer[103] [4]), .QN());
   DFF_X1 \o_buffer_reg[103][3]  (.D(n_123_707), .CK(n_120), .Q(
      \o_buffer[103] [3]), .QN());
   DFF_X1 \o_buffer_reg[103][2]  (.D(n_123_706), .CK(n_120), .Q(
      \o_buffer[103] [2]), .QN());
   DFF_X1 \o_buffer_reg[103][1]  (.D(n_123_705), .CK(n_120), .Q(
      \o_buffer[103] [1]), .QN());
   DFF_X1 \o_buffer_reg[103][0]  (.D(n_123_704), .CK(n_120), .Q(
      \o_buffer[103] [0]), .QN());
   DFF_X1 \o_buffer_reg[102][15]  (.D(n_123_703), .CK(n_120), .Q(
      \o_buffer[102] [15]), .QN());
   DFF_X1 \o_buffer_reg[102][14]  (.D(n_123_702), .CK(n_120), .Q(
      \o_buffer[102] [14]), .QN());
   DFF_X1 \o_buffer_reg[102][13]  (.D(n_123_701), .CK(n_120), .Q(
      \o_buffer[102] [13]), .QN());
   DFF_X1 \o_buffer_reg[102][12]  (.D(n_123_700), .CK(n_120), .Q(
      \o_buffer[102] [12]), .QN());
   DFF_X1 \o_buffer_reg[102][11]  (.D(n_123_699), .CK(n_120), .Q(
      \o_buffer[102] [11]), .QN());
   DFF_X1 \o_buffer_reg[102][10]  (.D(n_123_698), .CK(n_120), .Q(
      \o_buffer[102] [10]), .QN());
   DFF_X1 \o_buffer_reg[102][9]  (.D(n_123_697), .CK(n_120), .Q(
      \o_buffer[102] [9]), .QN());
   DFF_X1 \o_buffer_reg[102][8]  (.D(n_123_696), .CK(n_120), .Q(
      \o_buffer[102] [8]), .QN());
   DFF_X1 \o_buffer_reg[102][7]  (.D(n_123_695), .CK(n_120), .Q(
      \o_buffer[102] [7]), .QN());
   DFF_X1 \o_buffer_reg[102][6]  (.D(n_123_694), .CK(n_120), .Q(
      \o_buffer[102] [6]), .QN());
   DFF_X1 \o_buffer_reg[102][5]  (.D(n_123_693), .CK(n_120), .Q(
      \o_buffer[102] [5]), .QN());
   DFF_X1 \o_buffer_reg[102][4]  (.D(n_123_692), .CK(n_120), .Q(
      \o_buffer[102] [4]), .QN());
   DFF_X1 \o_buffer_reg[102][3]  (.D(n_123_691), .CK(n_120), .Q(
      \o_buffer[102] [3]), .QN());
   DFF_X1 \o_buffer_reg[102][2]  (.D(n_123_690), .CK(n_120), .Q(
      \o_buffer[102] [2]), .QN());
   DFF_X1 \o_buffer_reg[102][1]  (.D(n_123_689), .CK(n_120), .Q(
      \o_buffer[102] [1]), .QN());
   DFF_X1 \o_buffer_reg[102][0]  (.D(n_123_688), .CK(n_120), .Q(
      \o_buffer[102] [0]), .QN());
   DFF_X1 \o_buffer_reg[101][15]  (.D(n_123_687), .CK(n_120), .Q(
      \o_buffer[101] [15]), .QN());
   DFF_X1 \o_buffer_reg[101][14]  (.D(n_123_686), .CK(n_120), .Q(
      \o_buffer[101] [14]), .QN());
   DFF_X1 \o_buffer_reg[101][13]  (.D(n_123_685), .CK(n_120), .Q(
      \o_buffer[101] [13]), .QN());
   DFF_X1 \o_buffer_reg[101][12]  (.D(n_123_684), .CK(n_120), .Q(
      \o_buffer[101] [12]), .QN());
   DFF_X1 \o_buffer_reg[101][11]  (.D(n_123_683), .CK(n_120), .Q(
      \o_buffer[101] [11]), .QN());
   DFF_X1 \o_buffer_reg[101][10]  (.D(n_123_682), .CK(n_120), .Q(
      \o_buffer[101] [10]), .QN());
   DFF_X1 \o_buffer_reg[101][9]  (.D(n_123_681), .CK(n_120), .Q(
      \o_buffer[101] [9]), .QN());
   DFF_X1 \o_buffer_reg[101][8]  (.D(n_123_680), .CK(n_120), .Q(
      \o_buffer[101] [8]), .QN());
   DFF_X1 \o_buffer_reg[101][7]  (.D(n_123_679), .CK(n_120), .Q(
      \o_buffer[101] [7]), .QN());
   DFF_X1 \o_buffer_reg[101][6]  (.D(n_123_678), .CK(n_120), .Q(
      \o_buffer[101] [6]), .QN());
   DFF_X1 \o_buffer_reg[101][5]  (.D(n_123_677), .CK(n_120), .Q(
      \o_buffer[101] [5]), .QN());
   DFF_X1 \o_buffer_reg[101][4]  (.D(n_123_676), .CK(n_120), .Q(
      \o_buffer[101] [4]), .QN());
   DFF_X1 \o_buffer_reg[101][3]  (.D(n_123_675), .CK(n_120), .Q(
      \o_buffer[101] [3]), .QN());
   DFF_X1 \o_buffer_reg[101][2]  (.D(n_123_674), .CK(n_120), .Q(
      \o_buffer[101] [2]), .QN());
   DFF_X1 \o_buffer_reg[101][1]  (.D(n_123_673), .CK(n_120), .Q(
      \o_buffer[101] [1]), .QN());
   DFF_X1 \o_buffer_reg[101][0]  (.D(n_123_672), .CK(n_120), .Q(
      \o_buffer[101] [0]), .QN());
   DFF_X1 \o_buffer_reg[100][15]  (.D(n_123_671), .CK(n_120), .Q(
      \o_buffer[100] [15]), .QN());
   DFF_X1 \o_buffer_reg[100][14]  (.D(n_123_670), .CK(n_120), .Q(
      \o_buffer[100] [14]), .QN());
   DFF_X1 \o_buffer_reg[100][13]  (.D(n_123_669), .CK(n_120), .Q(
      \o_buffer[100] [13]), .QN());
   DFF_X1 \o_buffer_reg[100][12]  (.D(n_123_668), .CK(n_120), .Q(
      \o_buffer[100] [12]), .QN());
   DFF_X1 \o_buffer_reg[100][11]  (.D(n_123_667), .CK(n_120), .Q(
      \o_buffer[100] [11]), .QN());
   DFF_X1 \o_buffer_reg[100][10]  (.D(n_123_666), .CK(n_120), .Q(
      \o_buffer[100] [10]), .QN());
   DFF_X1 \o_buffer_reg[100][9]  (.D(n_123_665), .CK(n_120), .Q(
      \o_buffer[100] [9]), .QN());
   DFF_X1 \o_buffer_reg[100][8]  (.D(n_123_664), .CK(n_120), .Q(
      \o_buffer[100] [8]), .QN());
   DFF_X1 \o_buffer_reg[100][7]  (.D(n_123_663), .CK(n_120), .Q(
      \o_buffer[100] [7]), .QN());
   DFF_X1 \o_buffer_reg[100][6]  (.D(n_123_662), .CK(n_120), .Q(
      \o_buffer[100] [6]), .QN());
   DFF_X1 \o_buffer_reg[100][5]  (.D(n_123_661), .CK(n_120), .Q(
      \o_buffer[100] [5]), .QN());
   DFF_X1 \o_buffer_reg[100][4]  (.D(n_123_660), .CK(n_120), .Q(
      \o_buffer[100] [4]), .QN());
   DFF_X1 \o_buffer_reg[100][3]  (.D(n_123_659), .CK(n_120), .Q(
      \o_buffer[100] [3]), .QN());
   DFF_X1 \o_buffer_reg[100][2]  (.D(n_123_658), .CK(n_120), .Q(
      \o_buffer[100] [2]), .QN());
   DFF_X1 \o_buffer_reg[100][1]  (.D(n_123_657), .CK(n_120), .Q(
      \o_buffer[100] [1]), .QN());
   DFF_X1 \o_buffer_reg[100][0]  (.D(n_123_656), .CK(n_120), .Q(
      \o_buffer[100] [0]), .QN());
   DFF_X1 \o_buffer_reg[99][15]  (.D(n_123_655), .CK(n_120), .Q(
      \o_buffer[99] [15]), .QN());
   DFF_X1 \o_buffer_reg[99][14]  (.D(n_123_654), .CK(n_120), .Q(
      \o_buffer[99] [14]), .QN());
   DFF_X1 \o_buffer_reg[99][13]  (.D(n_123_653), .CK(n_120), .Q(
      \o_buffer[99] [13]), .QN());
   DFF_X1 \o_buffer_reg[99][12]  (.D(n_123_652), .CK(n_120), .Q(
      \o_buffer[99] [12]), .QN());
   DFF_X1 \o_buffer_reg[99][11]  (.D(n_123_651), .CK(n_120), .Q(
      \o_buffer[99] [11]), .QN());
   DFF_X1 \o_buffer_reg[99][10]  (.D(n_123_650), .CK(n_120), .Q(
      \o_buffer[99] [10]), .QN());
   DFF_X1 \o_buffer_reg[99][9]  (.D(n_123_649), .CK(n_120), .Q(\o_buffer[99] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][8]  (.D(n_123_648), .CK(n_120), .Q(\o_buffer[99] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][7]  (.D(n_123_647), .CK(n_120), .Q(\o_buffer[99] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][6]  (.D(n_123_646), .CK(n_120), .Q(\o_buffer[99] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][5]  (.D(n_123_645), .CK(n_120), .Q(\o_buffer[99] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][4]  (.D(n_123_644), .CK(n_120), .Q(\o_buffer[99] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][3]  (.D(n_123_643), .CK(n_120), .Q(\o_buffer[99] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][2]  (.D(n_123_642), .CK(n_120), .Q(\o_buffer[99] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][1]  (.D(n_123_641), .CK(n_120), .Q(\o_buffer[99] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[99][0]  (.D(n_123_640), .CK(n_120), .Q(\o_buffer[99] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][15]  (.D(n_123_639), .CK(n_120), .Q(
      \o_buffer[98] [15]), .QN());
   DFF_X1 \o_buffer_reg[98][14]  (.D(n_123_638), .CK(n_120), .Q(
      \o_buffer[98] [14]), .QN());
   DFF_X1 \o_buffer_reg[98][13]  (.D(n_123_637), .CK(n_120), .Q(
      \o_buffer[98] [13]), .QN());
   DFF_X1 \o_buffer_reg[98][12]  (.D(n_123_636), .CK(n_120), .Q(
      \o_buffer[98] [12]), .QN());
   DFF_X1 \o_buffer_reg[98][11]  (.D(n_123_635), .CK(n_120), .Q(
      \o_buffer[98] [11]), .QN());
   DFF_X1 \o_buffer_reg[98][10]  (.D(n_123_634), .CK(n_120), .Q(
      \o_buffer[98] [10]), .QN());
   DFF_X1 \o_buffer_reg[98][9]  (.D(n_123_633), .CK(n_120), .Q(\o_buffer[98] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][8]  (.D(n_123_632), .CK(n_120), .Q(\o_buffer[98] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][7]  (.D(n_123_631), .CK(n_120), .Q(\o_buffer[98] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][6]  (.D(n_123_630), .CK(n_120), .Q(\o_buffer[98] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][5]  (.D(n_123_629), .CK(n_120), .Q(\o_buffer[98] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][4]  (.D(n_123_628), .CK(n_120), .Q(\o_buffer[98] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][3]  (.D(n_123_627), .CK(n_120), .Q(\o_buffer[98] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][2]  (.D(n_123_626), .CK(n_120), .Q(\o_buffer[98] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][1]  (.D(n_123_625), .CK(n_120), .Q(\o_buffer[98] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[98][0]  (.D(n_123_624), .CK(n_120), .Q(\o_buffer[98] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][15]  (.D(n_123_623), .CK(n_120), .Q(
      \o_buffer[97] [15]), .QN());
   DFF_X1 \o_buffer_reg[97][14]  (.D(n_123_622), .CK(n_120), .Q(
      \o_buffer[97] [14]), .QN());
   DFF_X1 \o_buffer_reg[97][13]  (.D(n_123_621), .CK(n_120), .Q(
      \o_buffer[97] [13]), .QN());
   DFF_X1 \o_buffer_reg[97][12]  (.D(n_123_620), .CK(n_120), .Q(
      \o_buffer[97] [12]), .QN());
   DFF_X1 \o_buffer_reg[97][11]  (.D(n_123_619), .CK(n_120), .Q(
      \o_buffer[97] [11]), .QN());
   DFF_X1 \o_buffer_reg[97][10]  (.D(n_123_618), .CK(n_120), .Q(
      \o_buffer[97] [10]), .QN());
   DFF_X1 \o_buffer_reg[97][9]  (.D(n_123_617), .CK(n_120), .Q(\o_buffer[97] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][8]  (.D(n_123_616), .CK(n_120), .Q(\o_buffer[97] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][7]  (.D(n_123_615), .CK(n_120), .Q(\o_buffer[97] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][6]  (.D(n_123_614), .CK(n_120), .Q(\o_buffer[97] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][5]  (.D(n_123_613), .CK(n_120), .Q(\o_buffer[97] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][4]  (.D(n_123_612), .CK(n_120), .Q(\o_buffer[97] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][3]  (.D(n_123_611), .CK(n_120), .Q(\o_buffer[97] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][2]  (.D(n_123_610), .CK(n_120), .Q(\o_buffer[97] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][1]  (.D(n_123_609), .CK(n_120), .Q(\o_buffer[97] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[97][0]  (.D(n_123_608), .CK(n_120), .Q(\o_buffer[97] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][15]  (.D(n_123_607), .CK(n_120), .Q(
      \o_buffer[96] [15]), .QN());
   DFF_X1 \o_buffer_reg[96][14]  (.D(n_123_606), .CK(n_120), .Q(
      \o_buffer[96] [14]), .QN());
   DFF_X1 \o_buffer_reg[96][13]  (.D(n_123_605), .CK(n_120), .Q(
      \o_buffer[96] [13]), .QN());
   DFF_X1 \o_buffer_reg[96][12]  (.D(n_123_604), .CK(n_120), .Q(
      \o_buffer[96] [12]), .QN());
   DFF_X1 \o_buffer_reg[96][11]  (.D(n_123_603), .CK(n_120), .Q(
      \o_buffer[96] [11]), .QN());
   DFF_X1 \o_buffer_reg[96][10]  (.D(n_123_602), .CK(n_120), .Q(
      \o_buffer[96] [10]), .QN());
   DFF_X1 \o_buffer_reg[96][9]  (.D(n_123_601), .CK(n_120), .Q(\o_buffer[96] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][8]  (.D(n_123_600), .CK(n_120), .Q(\o_buffer[96] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][7]  (.D(n_123_599), .CK(n_120), .Q(\o_buffer[96] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][6]  (.D(n_123_598), .CK(n_120), .Q(\o_buffer[96] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][5]  (.D(n_123_597), .CK(n_120), .Q(\o_buffer[96] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][4]  (.D(n_123_596), .CK(n_120), .Q(\o_buffer[96] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][3]  (.D(n_123_595), .CK(n_120), .Q(\o_buffer[96] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][2]  (.D(n_123_594), .CK(n_120), .Q(\o_buffer[96] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][1]  (.D(n_123_593), .CK(n_120), .Q(\o_buffer[96] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[96][0]  (.D(n_123_592), .CK(n_120), .Q(\o_buffer[96] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][15]  (.D(n_123_591), .CK(n_120), .Q(
      \o_buffer[95] [15]), .QN());
   DFF_X1 \o_buffer_reg[95][14]  (.D(n_123_590), .CK(n_120), .Q(
      \o_buffer[95] [14]), .QN());
   DFF_X1 \o_buffer_reg[95][13]  (.D(n_123_589), .CK(n_120), .Q(
      \o_buffer[95] [13]), .QN());
   DFF_X1 \o_buffer_reg[95][12]  (.D(n_123_588), .CK(n_120), .Q(
      \o_buffer[95] [12]), .QN());
   DFF_X1 \o_buffer_reg[95][11]  (.D(n_123_587), .CK(n_120), .Q(
      \o_buffer[95] [11]), .QN());
   DFF_X1 \o_buffer_reg[95][10]  (.D(n_123_586), .CK(n_120), .Q(
      \o_buffer[95] [10]), .QN());
   DFF_X1 \o_buffer_reg[95][9]  (.D(n_123_585), .CK(n_120), .Q(\o_buffer[95] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][8]  (.D(n_123_584), .CK(n_120), .Q(\o_buffer[95] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][7]  (.D(n_123_583), .CK(n_120), .Q(\o_buffer[95] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][6]  (.D(n_123_582), .CK(n_120), .Q(\o_buffer[95] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][5]  (.D(n_123_581), .CK(n_120), .Q(\o_buffer[95] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][4]  (.D(n_123_580), .CK(n_120), .Q(\o_buffer[95] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][3]  (.D(n_123_579), .CK(n_120), .Q(\o_buffer[95] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][2]  (.D(n_123_578), .CK(n_120), .Q(\o_buffer[95] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][1]  (.D(n_123_577), .CK(n_120), .Q(\o_buffer[95] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[95][0]  (.D(n_123_576), .CK(n_120), .Q(\o_buffer[95] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][15]  (.D(n_123_575), .CK(n_120), .Q(
      \o_buffer[94] [15]), .QN());
   DFF_X1 \o_buffer_reg[94][14]  (.D(n_123_574), .CK(n_120), .Q(
      \o_buffer[94] [14]), .QN());
   DFF_X1 \o_buffer_reg[94][13]  (.D(n_123_573), .CK(n_120), .Q(
      \o_buffer[94] [13]), .QN());
   DFF_X1 \o_buffer_reg[94][12]  (.D(n_123_572), .CK(n_120), .Q(
      \o_buffer[94] [12]), .QN());
   DFF_X1 \o_buffer_reg[94][11]  (.D(n_123_571), .CK(n_120), .Q(
      \o_buffer[94] [11]), .QN());
   DFF_X1 \o_buffer_reg[94][10]  (.D(n_123_570), .CK(n_120), .Q(
      \o_buffer[94] [10]), .QN());
   DFF_X1 \o_buffer_reg[94][9]  (.D(n_123_569), .CK(n_120), .Q(\o_buffer[94] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][8]  (.D(n_123_568), .CK(n_120), .Q(\o_buffer[94] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][7]  (.D(n_123_567), .CK(n_120), .Q(\o_buffer[94] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][6]  (.D(n_123_566), .CK(n_120), .Q(\o_buffer[94] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][5]  (.D(n_123_565), .CK(n_120), .Q(\o_buffer[94] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][4]  (.D(n_123_564), .CK(n_120), .Q(\o_buffer[94] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][3]  (.D(n_123_563), .CK(n_120), .Q(\o_buffer[94] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][2]  (.D(n_123_562), .CK(n_120), .Q(\o_buffer[94] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][1]  (.D(n_123_561), .CK(n_120), .Q(\o_buffer[94] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[94][0]  (.D(n_123_560), .CK(n_120), .Q(\o_buffer[94] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][15]  (.D(n_123_559), .CK(n_120), .Q(
      \o_buffer[93] [15]), .QN());
   DFF_X1 \o_buffer_reg[93][14]  (.D(n_123_558), .CK(n_120), .Q(
      \o_buffer[93] [14]), .QN());
   DFF_X1 \o_buffer_reg[93][13]  (.D(n_123_557), .CK(n_120), .Q(
      \o_buffer[93] [13]), .QN());
   DFF_X1 \o_buffer_reg[93][12]  (.D(n_123_556), .CK(n_120), .Q(
      \o_buffer[93] [12]), .QN());
   DFF_X1 \o_buffer_reg[93][11]  (.D(n_123_555), .CK(n_120), .Q(
      \o_buffer[93] [11]), .QN());
   DFF_X1 \o_buffer_reg[93][10]  (.D(n_123_554), .CK(n_120), .Q(
      \o_buffer[93] [10]), .QN());
   DFF_X1 \o_buffer_reg[93][9]  (.D(n_123_553), .CK(n_120), .Q(\o_buffer[93] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][8]  (.D(n_123_552), .CK(n_120), .Q(\o_buffer[93] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][7]  (.D(n_123_551), .CK(n_120), .Q(\o_buffer[93] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][6]  (.D(n_123_550), .CK(n_120), .Q(\o_buffer[93] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][5]  (.D(n_123_549), .CK(n_120), .Q(\o_buffer[93] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][4]  (.D(n_123_548), .CK(n_120), .Q(\o_buffer[93] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][3]  (.D(n_123_547), .CK(n_120), .Q(\o_buffer[93] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][2]  (.D(n_123_546), .CK(n_120), .Q(\o_buffer[93] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][1]  (.D(n_123_545), .CK(n_120), .Q(\o_buffer[93] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[93][0]  (.D(n_123_544), .CK(n_120), .Q(\o_buffer[93] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][15]  (.D(n_123_543), .CK(n_120), .Q(
      \o_buffer[92] [15]), .QN());
   DFF_X1 \o_buffer_reg[92][14]  (.D(n_123_542), .CK(n_120), .Q(
      \o_buffer[92] [14]), .QN());
   DFF_X1 \o_buffer_reg[92][13]  (.D(n_123_541), .CK(n_120), .Q(
      \o_buffer[92] [13]), .QN());
   DFF_X1 \o_buffer_reg[92][12]  (.D(n_123_540), .CK(n_120), .Q(
      \o_buffer[92] [12]), .QN());
   DFF_X1 \o_buffer_reg[92][11]  (.D(n_123_539), .CK(n_120), .Q(
      \o_buffer[92] [11]), .QN());
   DFF_X1 \o_buffer_reg[92][10]  (.D(n_123_538), .CK(n_120), .Q(
      \o_buffer[92] [10]), .QN());
   DFF_X1 \o_buffer_reg[92][9]  (.D(n_123_537), .CK(n_120), .Q(\o_buffer[92] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][8]  (.D(n_123_536), .CK(n_120), .Q(\o_buffer[92] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][7]  (.D(n_123_535), .CK(n_120), .Q(\o_buffer[92] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][6]  (.D(n_123_534), .CK(n_120), .Q(\o_buffer[92] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][5]  (.D(n_123_533), .CK(n_120), .Q(\o_buffer[92] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][4]  (.D(n_123_532), .CK(n_120), .Q(\o_buffer[92] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][3]  (.D(n_123_531), .CK(n_120), .Q(\o_buffer[92] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][2]  (.D(n_123_530), .CK(n_120), .Q(\o_buffer[92] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][1]  (.D(n_123_529), .CK(n_120), .Q(\o_buffer[92] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[92][0]  (.D(n_123_528), .CK(n_120), .Q(\o_buffer[92] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][15]  (.D(n_123_527), .CK(n_120), .Q(
      \o_buffer[91] [15]), .QN());
   DFF_X1 \o_buffer_reg[91][14]  (.D(n_123_526), .CK(n_120), .Q(
      \o_buffer[91] [14]), .QN());
   DFF_X1 \o_buffer_reg[91][13]  (.D(n_123_525), .CK(n_120), .Q(
      \o_buffer[91] [13]), .QN());
   DFF_X1 \o_buffer_reg[91][12]  (.D(n_123_524), .CK(n_120), .Q(
      \o_buffer[91] [12]), .QN());
   DFF_X1 \o_buffer_reg[91][11]  (.D(n_123_523), .CK(n_120), .Q(
      \o_buffer[91] [11]), .QN());
   DFF_X1 \o_buffer_reg[91][10]  (.D(n_123_522), .CK(n_120), .Q(
      \o_buffer[91] [10]), .QN());
   DFF_X1 \o_buffer_reg[91][9]  (.D(n_123_521), .CK(n_120), .Q(\o_buffer[91] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][8]  (.D(n_123_520), .CK(n_120), .Q(\o_buffer[91] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][7]  (.D(n_123_519), .CK(n_120), .Q(\o_buffer[91] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][6]  (.D(n_123_518), .CK(n_120), .Q(\o_buffer[91] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][5]  (.D(n_123_517), .CK(n_120), .Q(\o_buffer[91] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][4]  (.D(n_123_516), .CK(n_120), .Q(\o_buffer[91] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][3]  (.D(n_123_515), .CK(n_120), .Q(\o_buffer[91] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][2]  (.D(n_123_514), .CK(n_120), .Q(\o_buffer[91] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][1]  (.D(n_123_513), .CK(n_120), .Q(\o_buffer[91] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[91][0]  (.D(n_123_512), .CK(n_120), .Q(\o_buffer[91] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][15]  (.D(n_123_511), .CK(n_120), .Q(
      \o_buffer[90] [15]), .QN());
   DFF_X1 \o_buffer_reg[90][14]  (.D(n_123_510), .CK(n_120), .Q(
      \o_buffer[90] [14]), .QN());
   DFF_X1 \o_buffer_reg[90][13]  (.D(n_123_509), .CK(n_120), .Q(
      \o_buffer[90] [13]), .QN());
   DFF_X1 \o_buffer_reg[90][12]  (.D(n_123_508), .CK(n_120), .Q(
      \o_buffer[90] [12]), .QN());
   DFF_X1 \o_buffer_reg[90][11]  (.D(n_123_507), .CK(n_120), .Q(
      \o_buffer[90] [11]), .QN());
   DFF_X1 \o_buffer_reg[90][10]  (.D(n_123_506), .CK(n_120), .Q(
      \o_buffer[90] [10]), .QN());
   DFF_X1 \o_buffer_reg[90][9]  (.D(n_123_505), .CK(n_120), .Q(\o_buffer[90] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][8]  (.D(n_123_504), .CK(n_120), .Q(\o_buffer[90] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][7]  (.D(n_123_503), .CK(n_120), .Q(\o_buffer[90] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][6]  (.D(n_123_502), .CK(n_120), .Q(\o_buffer[90] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][5]  (.D(n_123_501), .CK(n_120), .Q(\o_buffer[90] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][4]  (.D(n_123_500), .CK(n_120), .Q(\o_buffer[90] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][3]  (.D(n_123_499), .CK(n_120), .Q(\o_buffer[90] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][2]  (.D(n_123_498), .CK(n_120), .Q(\o_buffer[90] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][1]  (.D(n_123_497), .CK(n_120), .Q(\o_buffer[90] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[90][0]  (.D(n_123_496), .CK(n_120), .Q(\o_buffer[90] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][15]  (.D(n_123_495), .CK(n_120), .Q(
      \o_buffer[89] [15]), .QN());
   DFF_X1 \o_buffer_reg[89][14]  (.D(n_123_494), .CK(n_120), .Q(
      \o_buffer[89] [14]), .QN());
   DFF_X1 \o_buffer_reg[89][13]  (.D(n_123_493), .CK(n_120), .Q(
      \o_buffer[89] [13]), .QN());
   DFF_X1 \o_buffer_reg[89][12]  (.D(n_123_492), .CK(n_120), .Q(
      \o_buffer[89] [12]), .QN());
   DFF_X1 \o_buffer_reg[89][11]  (.D(n_123_491), .CK(n_120), .Q(
      \o_buffer[89] [11]), .QN());
   DFF_X1 \o_buffer_reg[89][10]  (.D(n_123_490), .CK(n_120), .Q(
      \o_buffer[89] [10]), .QN());
   DFF_X1 \o_buffer_reg[89][9]  (.D(n_123_489), .CK(n_120), .Q(\o_buffer[89] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][8]  (.D(n_123_488), .CK(n_120), .Q(\o_buffer[89] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][7]  (.D(n_123_487), .CK(n_120), .Q(\o_buffer[89] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][6]  (.D(n_123_486), .CK(n_120), .Q(\o_buffer[89] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][5]  (.D(n_123_485), .CK(n_120), .Q(\o_buffer[89] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][4]  (.D(n_123_484), .CK(n_120), .Q(\o_buffer[89] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][3]  (.D(n_123_483), .CK(n_120), .Q(\o_buffer[89] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][2]  (.D(n_123_482), .CK(n_120), .Q(\o_buffer[89] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][1]  (.D(n_123_481), .CK(n_120), .Q(\o_buffer[89] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[89][0]  (.D(n_123_480), .CK(n_120), .Q(\o_buffer[89] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][15]  (.D(n_123_479), .CK(n_120), .Q(
      \o_buffer[88] [15]), .QN());
   DFF_X1 \o_buffer_reg[88][14]  (.D(n_123_478), .CK(n_120), .Q(
      \o_buffer[88] [14]), .QN());
   DFF_X1 \o_buffer_reg[88][13]  (.D(n_123_477), .CK(n_120), .Q(
      \o_buffer[88] [13]), .QN());
   DFF_X1 \o_buffer_reg[88][12]  (.D(n_123_476), .CK(n_120), .Q(
      \o_buffer[88] [12]), .QN());
   DFF_X1 \o_buffer_reg[88][11]  (.D(n_123_475), .CK(n_120), .Q(
      \o_buffer[88] [11]), .QN());
   DFF_X1 \o_buffer_reg[88][10]  (.D(n_123_474), .CK(n_120), .Q(
      \o_buffer[88] [10]), .QN());
   DFF_X1 \o_buffer_reg[88][9]  (.D(n_123_473), .CK(n_120), .Q(\o_buffer[88] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][8]  (.D(n_123_472), .CK(n_120), .Q(\o_buffer[88] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][7]  (.D(n_123_471), .CK(n_120), .Q(\o_buffer[88] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][6]  (.D(n_123_470), .CK(n_120), .Q(\o_buffer[88] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][5]  (.D(n_123_469), .CK(n_120), .Q(\o_buffer[88] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][4]  (.D(n_123_468), .CK(n_120), .Q(\o_buffer[88] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][3]  (.D(n_123_467), .CK(n_120), .Q(\o_buffer[88] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][2]  (.D(n_123_466), .CK(n_120), .Q(\o_buffer[88] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][1]  (.D(n_123_465), .CK(n_120), .Q(\o_buffer[88] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[88][0]  (.D(n_123_464), .CK(n_120), .Q(\o_buffer[88] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][15]  (.D(n_123_463), .CK(n_120), .Q(
      \o_buffer[87] [15]), .QN());
   DFF_X1 \o_buffer_reg[87][14]  (.D(n_123_462), .CK(n_120), .Q(
      \o_buffer[87] [14]), .QN());
   DFF_X1 \o_buffer_reg[87][13]  (.D(n_123_461), .CK(n_120), .Q(
      \o_buffer[87] [13]), .QN());
   DFF_X1 \o_buffer_reg[87][12]  (.D(n_123_460), .CK(n_120), .Q(
      \o_buffer[87] [12]), .QN());
   DFF_X1 \o_buffer_reg[87][11]  (.D(n_123_459), .CK(n_120), .Q(
      \o_buffer[87] [11]), .QN());
   DFF_X1 \o_buffer_reg[87][10]  (.D(n_123_458), .CK(n_120), .Q(
      \o_buffer[87] [10]), .QN());
   DFF_X1 \o_buffer_reg[87][9]  (.D(n_123_457), .CK(n_120), .Q(\o_buffer[87] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][8]  (.D(n_123_456), .CK(n_120), .Q(\o_buffer[87] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][7]  (.D(n_123_455), .CK(n_120), .Q(\o_buffer[87] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][6]  (.D(n_123_454), .CK(n_120), .Q(\o_buffer[87] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][5]  (.D(n_123_453), .CK(n_120), .Q(\o_buffer[87] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][4]  (.D(n_123_452), .CK(n_120), .Q(\o_buffer[87] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][3]  (.D(n_123_451), .CK(n_120), .Q(\o_buffer[87] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][2]  (.D(n_123_450), .CK(n_120), .Q(\o_buffer[87] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][1]  (.D(n_123_449), .CK(n_120), .Q(\o_buffer[87] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[87][0]  (.D(n_123_448), .CK(n_120), .Q(\o_buffer[87] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][15]  (.D(n_123_447), .CK(n_120), .Q(
      \o_buffer[86] [15]), .QN());
   DFF_X1 \o_buffer_reg[86][14]  (.D(n_123_446), .CK(n_120), .Q(
      \o_buffer[86] [14]), .QN());
   DFF_X1 \o_buffer_reg[86][13]  (.D(n_123_445), .CK(n_120), .Q(
      \o_buffer[86] [13]), .QN());
   DFF_X1 \o_buffer_reg[86][12]  (.D(n_123_444), .CK(n_120), .Q(
      \o_buffer[86] [12]), .QN());
   DFF_X1 \o_buffer_reg[86][11]  (.D(n_123_443), .CK(n_120), .Q(
      \o_buffer[86] [11]), .QN());
   DFF_X1 \o_buffer_reg[86][10]  (.D(n_123_442), .CK(n_120), .Q(
      \o_buffer[86] [10]), .QN());
   DFF_X1 \o_buffer_reg[86][9]  (.D(n_123_441), .CK(n_120), .Q(\o_buffer[86] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][8]  (.D(n_123_440), .CK(n_120), .Q(\o_buffer[86] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][7]  (.D(n_123_439), .CK(n_120), .Q(\o_buffer[86] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][6]  (.D(n_123_438), .CK(n_120), .Q(\o_buffer[86] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][5]  (.D(n_123_437), .CK(n_120), .Q(\o_buffer[86] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][4]  (.D(n_123_436), .CK(n_120), .Q(\o_buffer[86] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][3]  (.D(n_123_435), .CK(n_120), .Q(\o_buffer[86] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][2]  (.D(n_123_434), .CK(n_120), .Q(\o_buffer[86] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][1]  (.D(n_123_433), .CK(n_120), .Q(\o_buffer[86] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[86][0]  (.D(n_123_432), .CK(n_120), .Q(\o_buffer[86] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][15]  (.D(n_123_431), .CK(n_120), .Q(
      \o_buffer[85] [15]), .QN());
   DFF_X1 \o_buffer_reg[85][14]  (.D(n_123_430), .CK(n_120), .Q(
      \o_buffer[85] [14]), .QN());
   DFF_X1 \o_buffer_reg[85][13]  (.D(n_123_429), .CK(n_120), .Q(
      \o_buffer[85] [13]), .QN());
   DFF_X1 \o_buffer_reg[85][12]  (.D(n_123_428), .CK(n_120), .Q(
      \o_buffer[85] [12]), .QN());
   DFF_X1 \o_buffer_reg[85][11]  (.D(n_123_427), .CK(n_120), .Q(
      \o_buffer[85] [11]), .QN());
   DFF_X1 \o_buffer_reg[85][10]  (.D(n_123_426), .CK(n_120), .Q(
      \o_buffer[85] [10]), .QN());
   DFF_X1 \o_buffer_reg[85][9]  (.D(n_123_425), .CK(n_120), .Q(\o_buffer[85] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][8]  (.D(n_123_424), .CK(n_120), .Q(\o_buffer[85] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][7]  (.D(n_123_423), .CK(n_120), .Q(\o_buffer[85] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][6]  (.D(n_123_422), .CK(n_120), .Q(\o_buffer[85] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][5]  (.D(n_123_421), .CK(n_120), .Q(\o_buffer[85] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][4]  (.D(n_123_420), .CK(n_120), .Q(\o_buffer[85] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][3]  (.D(n_123_419), .CK(n_120), .Q(\o_buffer[85] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][2]  (.D(n_123_418), .CK(n_120), .Q(\o_buffer[85] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][1]  (.D(n_123_417), .CK(n_120), .Q(\o_buffer[85] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[85][0]  (.D(n_123_416), .CK(n_120), .Q(\o_buffer[85] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][15]  (.D(n_123_415), .CK(n_120), .Q(
      \o_buffer[84] [15]), .QN());
   DFF_X1 \o_buffer_reg[84][14]  (.D(n_123_414), .CK(n_120), .Q(
      \o_buffer[84] [14]), .QN());
   DFF_X1 \o_buffer_reg[84][13]  (.D(n_123_413), .CK(n_120), .Q(
      \o_buffer[84] [13]), .QN());
   DFF_X1 \o_buffer_reg[84][12]  (.D(n_123_412), .CK(n_120), .Q(
      \o_buffer[84] [12]), .QN());
   DFF_X1 \o_buffer_reg[84][11]  (.D(n_123_411), .CK(n_120), .Q(
      \o_buffer[84] [11]), .QN());
   DFF_X1 \o_buffer_reg[84][10]  (.D(n_123_410), .CK(n_120), .Q(
      \o_buffer[84] [10]), .QN());
   DFF_X1 \o_buffer_reg[84][9]  (.D(n_123_409), .CK(n_120), .Q(\o_buffer[84] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][8]  (.D(n_123_408), .CK(n_120), .Q(\o_buffer[84] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][7]  (.D(n_123_407), .CK(n_120), .Q(\o_buffer[84] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][6]  (.D(n_123_406), .CK(n_120), .Q(\o_buffer[84] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][5]  (.D(n_123_405), .CK(n_120), .Q(\o_buffer[84] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][4]  (.D(n_123_404), .CK(n_120), .Q(\o_buffer[84] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][3]  (.D(n_123_403), .CK(n_120), .Q(\o_buffer[84] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][2]  (.D(n_123_402), .CK(n_120), .Q(\o_buffer[84] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][1]  (.D(n_123_401), .CK(n_120), .Q(\o_buffer[84] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[84][0]  (.D(n_123_400), .CK(n_120), .Q(\o_buffer[84] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][15]  (.D(n_123_399), .CK(n_120), .Q(
      \o_buffer[83] [15]), .QN());
   DFF_X1 \o_buffer_reg[83][14]  (.D(n_123_398), .CK(n_120), .Q(
      \o_buffer[83] [14]), .QN());
   DFF_X1 \o_buffer_reg[83][13]  (.D(n_123_397), .CK(n_120), .Q(
      \o_buffer[83] [13]), .QN());
   DFF_X1 \o_buffer_reg[83][12]  (.D(n_123_396), .CK(n_120), .Q(
      \o_buffer[83] [12]), .QN());
   DFF_X1 \o_buffer_reg[83][11]  (.D(n_123_395), .CK(n_120), .Q(
      \o_buffer[83] [11]), .QN());
   DFF_X1 \o_buffer_reg[83][10]  (.D(n_123_394), .CK(n_120), .Q(
      \o_buffer[83] [10]), .QN());
   DFF_X1 \o_buffer_reg[83][9]  (.D(n_123_393), .CK(n_120), .Q(\o_buffer[83] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][8]  (.D(n_123_392), .CK(n_120), .Q(\o_buffer[83] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][7]  (.D(n_123_391), .CK(n_120), .Q(\o_buffer[83] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][6]  (.D(n_123_390), .CK(n_120), .Q(\o_buffer[83] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][5]  (.D(n_123_389), .CK(n_120), .Q(\o_buffer[83] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][4]  (.D(n_123_388), .CK(n_120), .Q(\o_buffer[83] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][3]  (.D(n_123_387), .CK(n_120), .Q(\o_buffer[83] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][2]  (.D(n_123_386), .CK(n_120), .Q(\o_buffer[83] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][1]  (.D(n_123_385), .CK(n_120), .Q(\o_buffer[83] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[83][0]  (.D(n_123_384), .CK(n_120), .Q(\o_buffer[83] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][15]  (.D(n_123_383), .CK(n_120), .Q(
      \o_buffer[82] [15]), .QN());
   DFF_X1 \o_buffer_reg[82][14]  (.D(n_123_382), .CK(n_120), .Q(
      \o_buffer[82] [14]), .QN());
   DFF_X1 \o_buffer_reg[82][13]  (.D(n_123_381), .CK(n_120), .Q(
      \o_buffer[82] [13]), .QN());
   DFF_X1 \o_buffer_reg[82][12]  (.D(n_123_380), .CK(n_120), .Q(
      \o_buffer[82] [12]), .QN());
   DFF_X1 \o_buffer_reg[82][11]  (.D(n_123_379), .CK(n_120), .Q(
      \o_buffer[82] [11]), .QN());
   DFF_X1 \o_buffer_reg[82][10]  (.D(n_123_378), .CK(n_120), .Q(
      \o_buffer[82] [10]), .QN());
   DFF_X1 \o_buffer_reg[82][9]  (.D(n_123_377), .CK(n_120), .Q(\o_buffer[82] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][8]  (.D(n_123_376), .CK(n_120), .Q(\o_buffer[82] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][7]  (.D(n_123_375), .CK(n_120), .Q(\o_buffer[82] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][6]  (.D(n_123_374), .CK(n_120), .Q(\o_buffer[82] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][5]  (.D(n_123_373), .CK(n_120), .Q(\o_buffer[82] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][4]  (.D(n_123_372), .CK(n_120), .Q(\o_buffer[82] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][3]  (.D(n_123_371), .CK(n_120), .Q(\o_buffer[82] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][2]  (.D(n_123_370), .CK(n_120), .Q(\o_buffer[82] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][1]  (.D(n_123_369), .CK(n_120), .Q(\o_buffer[82] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[82][0]  (.D(n_123_368), .CK(n_120), .Q(\o_buffer[82] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][15]  (.D(n_123_367), .CK(n_120), .Q(
      \o_buffer[81] [15]), .QN());
   DFF_X1 \o_buffer_reg[81][14]  (.D(n_123_366), .CK(n_120), .Q(
      \o_buffer[81] [14]), .QN());
   DFF_X1 \o_buffer_reg[81][13]  (.D(n_123_365), .CK(n_120), .Q(
      \o_buffer[81] [13]), .QN());
   DFF_X1 \o_buffer_reg[81][12]  (.D(n_123_364), .CK(n_120), .Q(
      \o_buffer[81] [12]), .QN());
   DFF_X1 \o_buffer_reg[81][11]  (.D(n_123_363), .CK(n_120), .Q(
      \o_buffer[81] [11]), .QN());
   DFF_X1 \o_buffer_reg[81][10]  (.D(n_123_362), .CK(n_120), .Q(
      \o_buffer[81] [10]), .QN());
   DFF_X1 \o_buffer_reg[81][9]  (.D(n_123_361), .CK(n_120), .Q(\o_buffer[81] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][8]  (.D(n_123_360), .CK(n_120), .Q(\o_buffer[81] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][7]  (.D(n_123_359), .CK(n_120), .Q(\o_buffer[81] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][6]  (.D(n_123_358), .CK(n_120), .Q(\o_buffer[81] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][5]  (.D(n_123_357), .CK(n_120), .Q(\o_buffer[81] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][4]  (.D(n_123_356), .CK(n_120), .Q(\o_buffer[81] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][3]  (.D(n_123_355), .CK(n_120), .Q(\o_buffer[81] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][2]  (.D(n_123_354), .CK(n_120), .Q(\o_buffer[81] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][1]  (.D(n_123_353), .CK(n_120), .Q(\o_buffer[81] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[81][0]  (.D(n_123_352), .CK(n_120), .Q(\o_buffer[81] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][15]  (.D(n_123_351), .CK(n_120), .Q(
      \o_buffer[80] [15]), .QN());
   DFF_X1 \o_buffer_reg[80][14]  (.D(n_123_350), .CK(n_120), .Q(
      \o_buffer[80] [14]), .QN());
   DFF_X1 \o_buffer_reg[80][13]  (.D(n_123_349), .CK(n_120), .Q(
      \o_buffer[80] [13]), .QN());
   DFF_X1 \o_buffer_reg[80][12]  (.D(n_123_348), .CK(n_120), .Q(
      \o_buffer[80] [12]), .QN());
   DFF_X1 \o_buffer_reg[80][11]  (.D(n_123_347), .CK(n_120), .Q(
      \o_buffer[80] [11]), .QN());
   DFF_X1 \o_buffer_reg[80][10]  (.D(n_123_346), .CK(n_120), .Q(
      \o_buffer[80] [10]), .QN());
   DFF_X1 \o_buffer_reg[80][9]  (.D(n_123_345), .CK(n_120), .Q(\o_buffer[80] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][8]  (.D(n_123_344), .CK(n_120), .Q(\o_buffer[80] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][7]  (.D(n_123_343), .CK(n_120), .Q(\o_buffer[80] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][6]  (.D(n_123_342), .CK(n_120), .Q(\o_buffer[80] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][5]  (.D(n_123_341), .CK(n_120), .Q(\o_buffer[80] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][4]  (.D(n_123_340), .CK(n_120), .Q(\o_buffer[80] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][3]  (.D(n_123_339), .CK(n_120), .Q(\o_buffer[80] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][2]  (.D(n_123_338), .CK(n_120), .Q(\o_buffer[80] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][1]  (.D(n_123_337), .CK(n_120), .Q(\o_buffer[80] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[80][0]  (.D(n_123_336), .CK(n_120), .Q(\o_buffer[80] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][15]  (.D(n_123_335), .CK(n_120), .Q(
      \o_buffer[79] [15]), .QN());
   DFF_X1 \o_buffer_reg[79][14]  (.D(n_123_334), .CK(n_120), .Q(
      \o_buffer[79] [14]), .QN());
   DFF_X1 \o_buffer_reg[79][13]  (.D(n_123_333), .CK(n_120), .Q(
      \o_buffer[79] [13]), .QN());
   DFF_X1 \o_buffer_reg[79][12]  (.D(n_123_332), .CK(n_120), .Q(
      \o_buffer[79] [12]), .QN());
   DFF_X1 \o_buffer_reg[79][11]  (.D(n_123_331), .CK(n_120), .Q(
      \o_buffer[79] [11]), .QN());
   DFF_X1 \o_buffer_reg[79][10]  (.D(n_123_330), .CK(n_120), .Q(
      \o_buffer[79] [10]), .QN());
   DFF_X1 \o_buffer_reg[79][9]  (.D(n_123_329), .CK(n_120), .Q(\o_buffer[79] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][8]  (.D(n_123_328), .CK(n_120), .Q(\o_buffer[79] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][7]  (.D(n_123_327), .CK(n_120), .Q(\o_buffer[79] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][6]  (.D(n_123_326), .CK(n_120), .Q(\o_buffer[79] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][5]  (.D(n_123_325), .CK(n_120), .Q(\o_buffer[79] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][4]  (.D(n_123_324), .CK(n_120), .Q(\o_buffer[79] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][3]  (.D(n_123_323), .CK(n_120), .Q(\o_buffer[79] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][2]  (.D(n_123_322), .CK(n_120), .Q(\o_buffer[79] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][1]  (.D(n_123_321), .CK(n_120), .Q(\o_buffer[79] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[79][0]  (.D(n_123_320), .CK(n_120), .Q(\o_buffer[79] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][15]  (.D(n_123_319), .CK(n_120), .Q(
      \o_buffer[78] [15]), .QN());
   DFF_X1 \o_buffer_reg[78][14]  (.D(n_123_318), .CK(n_120), .Q(
      \o_buffer[78] [14]), .QN());
   DFF_X1 \o_buffer_reg[78][13]  (.D(n_123_317), .CK(n_120), .Q(
      \o_buffer[78] [13]), .QN());
   DFF_X1 \o_buffer_reg[78][12]  (.D(n_123_316), .CK(n_120), .Q(
      \o_buffer[78] [12]), .QN());
   DFF_X1 \o_buffer_reg[78][11]  (.D(n_123_315), .CK(n_120), .Q(
      \o_buffer[78] [11]), .QN());
   DFF_X1 \o_buffer_reg[78][10]  (.D(n_123_314), .CK(n_120), .Q(
      \o_buffer[78] [10]), .QN());
   DFF_X1 \o_buffer_reg[78][9]  (.D(n_123_313), .CK(n_120), .Q(\o_buffer[78] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][8]  (.D(n_123_312), .CK(n_120), .Q(\o_buffer[78] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][7]  (.D(n_123_311), .CK(n_120), .Q(\o_buffer[78] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][6]  (.D(n_123_310), .CK(n_120), .Q(\o_buffer[78] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][5]  (.D(n_123_309), .CK(n_120), .Q(\o_buffer[78] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][4]  (.D(n_123_308), .CK(n_120), .Q(\o_buffer[78] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][3]  (.D(n_123_307), .CK(n_120), .Q(\o_buffer[78] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][2]  (.D(n_123_306), .CK(n_120), .Q(\o_buffer[78] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][1]  (.D(n_123_305), .CK(n_120), .Q(\o_buffer[78] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[78][0]  (.D(n_123_304), .CK(n_120), .Q(\o_buffer[78] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][15]  (.D(n_123_303), .CK(n_120), .Q(
      \o_buffer[77] [15]), .QN());
   DFF_X1 \o_buffer_reg[77][14]  (.D(n_123_302), .CK(n_120), .Q(
      \o_buffer[77] [14]), .QN());
   DFF_X1 \o_buffer_reg[77][13]  (.D(n_123_301), .CK(n_120), .Q(
      \o_buffer[77] [13]), .QN());
   DFF_X1 \o_buffer_reg[77][12]  (.D(n_123_300), .CK(n_120), .Q(
      \o_buffer[77] [12]), .QN());
   DFF_X1 \o_buffer_reg[77][11]  (.D(n_123_299), .CK(n_120), .Q(
      \o_buffer[77] [11]), .QN());
   DFF_X1 \o_buffer_reg[77][10]  (.D(n_123_298), .CK(n_120), .Q(
      \o_buffer[77] [10]), .QN());
   DFF_X1 \o_buffer_reg[77][9]  (.D(n_123_297), .CK(n_120), .Q(\o_buffer[77] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][8]  (.D(n_123_296), .CK(n_120), .Q(\o_buffer[77] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][7]  (.D(n_123_295), .CK(n_120), .Q(\o_buffer[77] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][6]  (.D(n_123_294), .CK(n_120), .Q(\o_buffer[77] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][5]  (.D(n_123_293), .CK(n_120), .Q(\o_buffer[77] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][4]  (.D(n_123_292), .CK(n_120), .Q(\o_buffer[77] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][3]  (.D(n_123_291), .CK(n_120), .Q(\o_buffer[77] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][2]  (.D(n_123_290), .CK(n_120), .Q(\o_buffer[77] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][1]  (.D(n_123_289), .CK(n_120), .Q(\o_buffer[77] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[77][0]  (.D(n_123_288), .CK(n_120), .Q(\o_buffer[77] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][15]  (.D(n_123_287), .CK(n_120), .Q(
      \o_buffer[76] [15]), .QN());
   DFF_X1 \o_buffer_reg[76][14]  (.D(n_123_286), .CK(n_120), .Q(
      \o_buffer[76] [14]), .QN());
   DFF_X1 \o_buffer_reg[76][13]  (.D(n_123_285), .CK(n_120), .Q(
      \o_buffer[76] [13]), .QN());
   DFF_X1 \o_buffer_reg[76][12]  (.D(n_123_284), .CK(n_120), .Q(
      \o_buffer[76] [12]), .QN());
   DFF_X1 \o_buffer_reg[76][11]  (.D(n_123_283), .CK(n_120), .Q(
      \o_buffer[76] [11]), .QN());
   DFF_X1 \o_buffer_reg[76][10]  (.D(n_123_282), .CK(n_120), .Q(
      \o_buffer[76] [10]), .QN());
   DFF_X1 \o_buffer_reg[76][9]  (.D(n_123_281), .CK(n_120), .Q(\o_buffer[76] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][8]  (.D(n_123_280), .CK(n_120), .Q(\o_buffer[76] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][7]  (.D(n_123_279), .CK(n_120), .Q(\o_buffer[76] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][6]  (.D(n_123_278), .CK(n_120), .Q(\o_buffer[76] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][5]  (.D(n_123_277), .CK(n_120), .Q(\o_buffer[76] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][4]  (.D(n_123_276), .CK(n_120), .Q(\o_buffer[76] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][3]  (.D(n_123_275), .CK(n_120), .Q(\o_buffer[76] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][2]  (.D(n_123_274), .CK(n_120), .Q(\o_buffer[76] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][1]  (.D(n_123_273), .CK(n_120), .Q(\o_buffer[76] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[76][0]  (.D(n_123_272), .CK(n_120), .Q(\o_buffer[76] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][15]  (.D(n_123_271), .CK(n_120), .Q(
      \o_buffer[75] [15]), .QN());
   DFF_X1 \o_buffer_reg[75][14]  (.D(n_123_270), .CK(n_120), .Q(
      \o_buffer[75] [14]), .QN());
   DFF_X1 \o_buffer_reg[75][13]  (.D(n_123_269), .CK(n_120), .Q(
      \o_buffer[75] [13]), .QN());
   DFF_X1 \o_buffer_reg[75][12]  (.D(n_123_268), .CK(n_120), .Q(
      \o_buffer[75] [12]), .QN());
   DFF_X1 \o_buffer_reg[75][11]  (.D(n_123_267), .CK(n_120), .Q(
      \o_buffer[75] [11]), .QN());
   DFF_X1 \o_buffer_reg[75][10]  (.D(n_123_266), .CK(n_120), .Q(
      \o_buffer[75] [10]), .QN());
   DFF_X1 \o_buffer_reg[75][9]  (.D(n_123_265), .CK(n_120), .Q(\o_buffer[75] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][8]  (.D(n_123_264), .CK(n_120), .Q(\o_buffer[75] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][7]  (.D(n_123_263), .CK(n_120), .Q(\o_buffer[75] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][6]  (.D(n_123_262), .CK(n_120), .Q(\o_buffer[75] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][5]  (.D(n_123_261), .CK(n_120), .Q(\o_buffer[75] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][4]  (.D(n_123_260), .CK(n_120), .Q(\o_buffer[75] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][3]  (.D(n_123_259), .CK(n_120), .Q(\o_buffer[75] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][2]  (.D(n_123_258), .CK(n_120), .Q(\o_buffer[75] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][1]  (.D(n_123_257), .CK(n_120), .Q(\o_buffer[75] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[75][0]  (.D(n_123_256), .CK(n_120), .Q(\o_buffer[75] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][15]  (.D(n_123_255), .CK(n_120), .Q(
      \o_buffer[74] [15]), .QN());
   DFF_X1 \o_buffer_reg[74][14]  (.D(n_123_254), .CK(n_120), .Q(
      \o_buffer[74] [14]), .QN());
   DFF_X1 \o_buffer_reg[74][13]  (.D(n_123_253), .CK(n_120), .Q(
      \o_buffer[74] [13]), .QN());
   DFF_X1 \o_buffer_reg[74][12]  (.D(n_123_252), .CK(n_120), .Q(
      \o_buffer[74] [12]), .QN());
   DFF_X1 \o_buffer_reg[74][11]  (.D(n_123_251), .CK(n_120), .Q(
      \o_buffer[74] [11]), .QN());
   DFF_X1 \o_buffer_reg[74][10]  (.D(n_123_250), .CK(n_120), .Q(
      \o_buffer[74] [10]), .QN());
   DFF_X1 \o_buffer_reg[74][9]  (.D(n_123_249), .CK(n_120), .Q(\o_buffer[74] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][8]  (.D(n_123_248), .CK(n_120), .Q(\o_buffer[74] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][7]  (.D(n_123_247), .CK(n_120), .Q(\o_buffer[74] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][6]  (.D(n_123_246), .CK(n_120), .Q(\o_buffer[74] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][5]  (.D(n_123_245), .CK(n_120), .Q(\o_buffer[74] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][4]  (.D(n_123_244), .CK(n_120), .Q(\o_buffer[74] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][3]  (.D(n_123_243), .CK(n_120), .Q(\o_buffer[74] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][2]  (.D(n_123_242), .CK(n_120), .Q(\o_buffer[74] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][1]  (.D(n_123_241), .CK(n_120), .Q(\o_buffer[74] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[74][0]  (.D(n_123_240), .CK(n_120), .Q(\o_buffer[74] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][15]  (.D(n_123_239), .CK(n_120), .Q(
      \o_buffer[73] [15]), .QN());
   DFF_X1 \o_buffer_reg[73][14]  (.D(n_123_238), .CK(n_120), .Q(
      \o_buffer[73] [14]), .QN());
   DFF_X1 \o_buffer_reg[73][13]  (.D(n_123_237), .CK(n_120), .Q(
      \o_buffer[73] [13]), .QN());
   DFF_X1 \o_buffer_reg[73][12]  (.D(n_123_236), .CK(n_120), .Q(
      \o_buffer[73] [12]), .QN());
   DFF_X1 \o_buffer_reg[73][11]  (.D(n_123_235), .CK(n_120), .Q(
      \o_buffer[73] [11]), .QN());
   DFF_X1 \o_buffer_reg[73][10]  (.D(n_123_234), .CK(n_120), .Q(
      \o_buffer[73] [10]), .QN());
   DFF_X1 \o_buffer_reg[73][9]  (.D(n_123_233), .CK(n_120), .Q(\o_buffer[73] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][8]  (.D(n_123_232), .CK(n_120), .Q(\o_buffer[73] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][7]  (.D(n_123_231), .CK(n_120), .Q(\o_buffer[73] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][6]  (.D(n_123_230), .CK(n_120), .Q(\o_buffer[73] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][5]  (.D(n_123_229), .CK(n_120), .Q(\o_buffer[73] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][4]  (.D(n_123_228), .CK(n_120), .Q(\o_buffer[73] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][3]  (.D(n_123_227), .CK(n_120), .Q(\o_buffer[73] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][2]  (.D(n_123_226), .CK(n_120), .Q(\o_buffer[73] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][1]  (.D(n_123_225), .CK(n_120), .Q(\o_buffer[73] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[73][0]  (.D(n_123_224), .CK(n_120), .Q(\o_buffer[73] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][15]  (.D(n_123_223), .CK(n_120), .Q(
      \o_buffer[72] [15]), .QN());
   DFF_X1 \o_buffer_reg[72][14]  (.D(n_123_222), .CK(n_120), .Q(
      \o_buffer[72] [14]), .QN());
   DFF_X1 \o_buffer_reg[72][13]  (.D(n_123_221), .CK(n_120), .Q(
      \o_buffer[72] [13]), .QN());
   DFF_X1 \o_buffer_reg[72][12]  (.D(n_123_220), .CK(n_120), .Q(
      \o_buffer[72] [12]), .QN());
   DFF_X1 \o_buffer_reg[72][11]  (.D(n_123_219), .CK(n_120), .Q(
      \o_buffer[72] [11]), .QN());
   DFF_X1 \o_buffer_reg[72][10]  (.D(n_123_218), .CK(n_120), .Q(
      \o_buffer[72] [10]), .QN());
   DFF_X1 \o_buffer_reg[72][9]  (.D(n_123_217), .CK(n_120), .Q(\o_buffer[72] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][8]  (.D(n_123_216), .CK(n_120), .Q(\o_buffer[72] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][7]  (.D(n_123_215), .CK(n_120), .Q(\o_buffer[72] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][6]  (.D(n_123_214), .CK(n_120), .Q(\o_buffer[72] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][5]  (.D(n_123_213), .CK(n_120), .Q(\o_buffer[72] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][4]  (.D(n_123_212), .CK(n_120), .Q(\o_buffer[72] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][3]  (.D(n_123_211), .CK(n_120), .Q(\o_buffer[72] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][2]  (.D(n_123_210), .CK(n_120), .Q(\o_buffer[72] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][1]  (.D(n_123_209), .CK(n_120), .Q(\o_buffer[72] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[72][0]  (.D(n_123_208), .CK(n_120), .Q(\o_buffer[72] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][15]  (.D(n_123_207), .CK(n_120), .Q(
      \o_buffer[71] [15]), .QN());
   DFF_X1 \o_buffer_reg[71][14]  (.D(n_123_206), .CK(n_120), .Q(
      \o_buffer[71] [14]), .QN());
   DFF_X1 \o_buffer_reg[71][13]  (.D(n_123_205), .CK(n_120), .Q(
      \o_buffer[71] [13]), .QN());
   DFF_X1 \o_buffer_reg[71][12]  (.D(n_123_204), .CK(n_120), .Q(
      \o_buffer[71] [12]), .QN());
   DFF_X1 \o_buffer_reg[71][11]  (.D(n_123_203), .CK(n_120), .Q(
      \o_buffer[71] [11]), .QN());
   DFF_X1 \o_buffer_reg[71][10]  (.D(n_123_202), .CK(n_120), .Q(
      \o_buffer[71] [10]), .QN());
   DFF_X1 \o_buffer_reg[71][9]  (.D(n_123_201), .CK(n_120), .Q(\o_buffer[71] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][8]  (.D(n_123_200), .CK(n_120), .Q(\o_buffer[71] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][7]  (.D(n_123_199), .CK(n_120), .Q(\o_buffer[71] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][6]  (.D(n_123_198), .CK(n_120), .Q(\o_buffer[71] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][5]  (.D(n_123_197), .CK(n_120), .Q(\o_buffer[71] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][4]  (.D(n_123_196), .CK(n_120), .Q(\o_buffer[71] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][3]  (.D(n_123_195), .CK(n_120), .Q(\o_buffer[71] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][2]  (.D(n_123_194), .CK(n_120), .Q(\o_buffer[71] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][1]  (.D(n_123_193), .CK(n_120), .Q(\o_buffer[71] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[71][0]  (.D(n_123_192), .CK(n_120), .Q(\o_buffer[71] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][15]  (.D(n_123_191), .CK(n_120), .Q(
      \o_buffer[70] [15]), .QN());
   DFF_X1 \o_buffer_reg[70][14]  (.D(n_123_190), .CK(n_120), .Q(
      \o_buffer[70] [14]), .QN());
   DFF_X1 \o_buffer_reg[70][13]  (.D(n_123_189), .CK(n_120), .Q(
      \o_buffer[70] [13]), .QN());
   DFF_X1 \o_buffer_reg[70][12]  (.D(n_123_188), .CK(n_120), .Q(
      \o_buffer[70] [12]), .QN());
   DFF_X1 \o_buffer_reg[70][11]  (.D(n_123_187), .CK(n_120), .Q(
      \o_buffer[70] [11]), .QN());
   DFF_X1 \o_buffer_reg[70][10]  (.D(n_123_186), .CK(n_120), .Q(
      \o_buffer[70] [10]), .QN());
   DFF_X1 \o_buffer_reg[70][9]  (.D(n_123_185), .CK(n_120), .Q(\o_buffer[70] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][8]  (.D(n_123_184), .CK(n_120), .Q(\o_buffer[70] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][7]  (.D(n_123_183), .CK(n_120), .Q(\o_buffer[70] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][6]  (.D(n_123_182), .CK(n_120), .Q(\o_buffer[70] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][5]  (.D(n_123_181), .CK(n_120), .Q(\o_buffer[70] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][4]  (.D(n_123_180), .CK(n_120), .Q(\o_buffer[70] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][3]  (.D(n_123_179), .CK(n_120), .Q(\o_buffer[70] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][2]  (.D(n_123_178), .CK(n_120), .Q(\o_buffer[70] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][1]  (.D(n_123_177), .CK(n_120), .Q(\o_buffer[70] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[70][0]  (.D(n_123_176), .CK(n_120), .Q(\o_buffer[70] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][15]  (.D(n_123_175), .CK(n_120), .Q(
      \o_buffer[69] [15]), .QN());
   DFF_X1 \o_buffer_reg[69][14]  (.D(n_123_174), .CK(n_120), .Q(
      \o_buffer[69] [14]), .QN());
   DFF_X1 \o_buffer_reg[69][13]  (.D(n_123_173), .CK(n_120), .Q(
      \o_buffer[69] [13]), .QN());
   DFF_X1 \o_buffer_reg[69][12]  (.D(n_123_172), .CK(n_120), .Q(
      \o_buffer[69] [12]), .QN());
   DFF_X1 \o_buffer_reg[69][11]  (.D(n_123_171), .CK(n_120), .Q(
      \o_buffer[69] [11]), .QN());
   DFF_X1 \o_buffer_reg[69][10]  (.D(n_123_170), .CK(n_120), .Q(
      \o_buffer[69] [10]), .QN());
   DFF_X1 \o_buffer_reg[69][9]  (.D(n_123_169), .CK(n_120), .Q(\o_buffer[69] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][8]  (.D(n_123_168), .CK(n_120), .Q(\o_buffer[69] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][7]  (.D(n_123_167), .CK(n_120), .Q(\o_buffer[69] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][6]  (.D(n_123_166), .CK(n_120), .Q(\o_buffer[69] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][5]  (.D(n_123_165), .CK(n_120), .Q(\o_buffer[69] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][4]  (.D(n_123_164), .CK(n_120), .Q(\o_buffer[69] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][3]  (.D(n_123_163), .CK(n_120), .Q(\o_buffer[69] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][2]  (.D(n_123_162), .CK(n_120), .Q(\o_buffer[69] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][1]  (.D(n_123_161), .CK(n_120), .Q(\o_buffer[69] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[69][0]  (.D(n_123_160), .CK(n_120), .Q(\o_buffer[69] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][15]  (.D(n_123_159), .CK(n_120), .Q(
      \o_buffer[68] [15]), .QN());
   DFF_X1 \o_buffer_reg[68][14]  (.D(n_123_158), .CK(n_120), .Q(
      \o_buffer[68] [14]), .QN());
   DFF_X1 \o_buffer_reg[68][13]  (.D(n_123_157), .CK(n_120), .Q(
      \o_buffer[68] [13]), .QN());
   DFF_X1 \o_buffer_reg[68][12]  (.D(n_123_156), .CK(n_120), .Q(
      \o_buffer[68] [12]), .QN());
   DFF_X1 \o_buffer_reg[68][11]  (.D(n_123_155), .CK(n_120), .Q(
      \o_buffer[68] [11]), .QN());
   DFF_X1 \o_buffer_reg[68][10]  (.D(n_123_154), .CK(n_120), .Q(
      \o_buffer[68] [10]), .QN());
   DFF_X1 \o_buffer_reg[68][9]  (.D(n_123_153), .CK(n_120), .Q(\o_buffer[68] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][8]  (.D(n_123_152), .CK(n_120), .Q(\o_buffer[68] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][7]  (.D(n_123_151), .CK(n_120), .Q(\o_buffer[68] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][6]  (.D(n_123_150), .CK(n_120), .Q(\o_buffer[68] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][5]  (.D(n_123_149), .CK(n_120), .Q(\o_buffer[68] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][4]  (.D(n_123_148), .CK(n_120), .Q(\o_buffer[68] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][3]  (.D(n_123_147), .CK(n_120), .Q(\o_buffer[68] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][2]  (.D(n_123_146), .CK(n_120), .Q(\o_buffer[68] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][1]  (.D(n_123_145), .CK(n_120), .Q(\o_buffer[68] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[68][0]  (.D(n_123_144), .CK(n_120), .Q(\o_buffer[68] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][15]  (.D(n_123_143), .CK(n_120), .Q(
      \o_buffer[67] [15]), .QN());
   DFF_X1 \o_buffer_reg[67][14]  (.D(n_123_142), .CK(n_120), .Q(
      \o_buffer[67] [14]), .QN());
   DFF_X1 \o_buffer_reg[67][13]  (.D(n_123_141), .CK(n_120), .Q(
      \o_buffer[67] [13]), .QN());
   DFF_X1 \o_buffer_reg[67][12]  (.D(n_123_140), .CK(n_120), .Q(
      \o_buffer[67] [12]), .QN());
   DFF_X1 \o_buffer_reg[67][11]  (.D(n_123_139), .CK(n_120), .Q(
      \o_buffer[67] [11]), .QN());
   DFF_X1 \o_buffer_reg[67][10]  (.D(n_123_138), .CK(n_120), .Q(
      \o_buffer[67] [10]), .QN());
   DFF_X1 \o_buffer_reg[67][9]  (.D(n_123_137), .CK(n_120), .Q(\o_buffer[67] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][8]  (.D(n_123_136), .CK(n_120), .Q(\o_buffer[67] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][7]  (.D(n_123_135), .CK(n_120), .Q(\o_buffer[67] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][6]  (.D(n_123_134), .CK(n_120), .Q(\o_buffer[67] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][5]  (.D(n_123_133), .CK(n_120), .Q(\o_buffer[67] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][4]  (.D(n_123_132), .CK(n_120), .Q(\o_buffer[67] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][3]  (.D(n_123_131), .CK(n_120), .Q(\o_buffer[67] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][2]  (.D(n_123_130), .CK(n_120), .Q(\o_buffer[67] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][1]  (.D(n_123_129), .CK(n_120), .Q(\o_buffer[67] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[67][0]  (.D(n_123_128), .CK(n_120), .Q(\o_buffer[67] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][15]  (.D(n_123_127), .CK(n_120), .Q(
      \o_buffer[66] [15]), .QN());
   DFF_X1 \o_buffer_reg[66][14]  (.D(n_123_126), .CK(n_120), .Q(
      \o_buffer[66] [14]), .QN());
   DFF_X1 \o_buffer_reg[66][13]  (.D(n_123_125), .CK(n_120), .Q(
      \o_buffer[66] [13]), .QN());
   DFF_X1 \o_buffer_reg[66][12]  (.D(n_123_124), .CK(n_120), .Q(
      \o_buffer[66] [12]), .QN());
   DFF_X1 \o_buffer_reg[66][11]  (.D(n_123_123), .CK(n_120), .Q(
      \o_buffer[66] [11]), .QN());
   DFF_X1 \o_buffer_reg[66][10]  (.D(n_123_122), .CK(n_120), .Q(
      \o_buffer[66] [10]), .QN());
   DFF_X1 \o_buffer_reg[66][9]  (.D(n_123_121), .CK(n_120), .Q(\o_buffer[66] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][8]  (.D(n_123_120), .CK(n_120), .Q(\o_buffer[66] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][7]  (.D(n_123_119), .CK(n_120), .Q(\o_buffer[66] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][6]  (.D(n_123_118), .CK(n_120), .Q(\o_buffer[66] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][5]  (.D(n_123_117), .CK(n_120), .Q(\o_buffer[66] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][4]  (.D(n_123_116), .CK(n_120), .Q(\o_buffer[66] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][3]  (.D(n_123_115), .CK(n_120), .Q(\o_buffer[66] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][2]  (.D(n_123_114), .CK(n_120), .Q(\o_buffer[66] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][1]  (.D(n_123_113), .CK(n_120), .Q(\o_buffer[66] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[66][0]  (.D(n_123_112), .CK(n_120), .Q(\o_buffer[66] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][15]  (.D(n_123_111), .CK(n_120), .Q(
      \o_buffer[65] [15]), .QN());
   DFF_X1 \o_buffer_reg[65][14]  (.D(n_123_110), .CK(n_120), .Q(
      \o_buffer[65] [14]), .QN());
   DFF_X1 \o_buffer_reg[65][13]  (.D(n_123_109), .CK(n_120), .Q(
      \o_buffer[65] [13]), .QN());
   DFF_X1 \o_buffer_reg[65][12]  (.D(n_123_108), .CK(n_120), .Q(
      \o_buffer[65] [12]), .QN());
   DFF_X1 \o_buffer_reg[65][11]  (.D(n_123_107), .CK(n_120), .Q(
      \o_buffer[65] [11]), .QN());
   DFF_X1 \o_buffer_reg[65][10]  (.D(n_123_106), .CK(n_120), .Q(
      \o_buffer[65] [10]), .QN());
   DFF_X1 \o_buffer_reg[65][9]  (.D(n_123_105), .CK(n_120), .Q(\o_buffer[65] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][8]  (.D(n_123_104), .CK(n_120), .Q(\o_buffer[65] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][7]  (.D(n_123_103), .CK(n_120), .Q(\o_buffer[65] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][6]  (.D(n_123_102), .CK(n_120), .Q(\o_buffer[65] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][5]  (.D(n_123_101), .CK(n_120), .Q(\o_buffer[65] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][4]  (.D(n_123_100), .CK(n_120), .Q(\o_buffer[65] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][3]  (.D(n_123_99), .CK(n_120), .Q(\o_buffer[65] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][2]  (.D(n_123_98), .CK(n_120), .Q(\o_buffer[65] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][1]  (.D(n_123_97), .CK(n_120), .Q(\o_buffer[65] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[65][0]  (.D(n_123_96), .CK(n_120), .Q(\o_buffer[65] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][15]  (.D(n_123_95), .CK(n_120), .Q(
      \o_buffer[64] [15]), .QN());
   DFF_X1 \o_buffer_reg[64][14]  (.D(n_123_94), .CK(n_120), .Q(
      \o_buffer[64] [14]), .QN());
   DFF_X1 \o_buffer_reg[64][13]  (.D(n_123_93), .CK(n_120), .Q(
      \o_buffer[64] [13]), .QN());
   DFF_X1 \o_buffer_reg[64][12]  (.D(n_123_92), .CK(n_120), .Q(
      \o_buffer[64] [12]), .QN());
   DFF_X1 \o_buffer_reg[64][11]  (.D(n_123_91), .CK(n_120), .Q(
      \o_buffer[64] [11]), .QN());
   DFF_X1 \o_buffer_reg[64][10]  (.D(n_123_90), .CK(n_120), .Q(
      \o_buffer[64] [10]), .QN());
   DFF_X1 \o_buffer_reg[64][9]  (.D(n_123_89), .CK(n_120), .Q(\o_buffer[64] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][8]  (.D(n_123_88), .CK(n_120), .Q(\o_buffer[64] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][7]  (.D(n_123_87), .CK(n_120), .Q(\o_buffer[64] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][6]  (.D(n_123_86), .CK(n_120), .Q(\o_buffer[64] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][5]  (.D(n_123_85), .CK(n_120), .Q(\o_buffer[64] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][4]  (.D(n_123_84), .CK(n_120), .Q(\o_buffer[64] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][3]  (.D(n_123_83), .CK(n_120), .Q(\o_buffer[64] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][2]  (.D(n_123_82), .CK(n_120), .Q(\o_buffer[64] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][1]  (.D(n_123_81), .CK(n_120), .Q(\o_buffer[64] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[64][0]  (.D(n_123_80), .CK(n_120), .Q(\o_buffer[64] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][15]  (.D(n_123_79), .CK(n_120), .Q(
      \o_buffer[63] [15]), .QN());
   DFF_X1 \o_buffer_reg[63][14]  (.D(n_123_78), .CK(n_120), .Q(
      \o_buffer[63] [14]), .QN());
   DFF_X1 \o_buffer_reg[63][13]  (.D(n_123_77), .CK(n_120), .Q(
      \o_buffer[63] [13]), .QN());
   DFF_X1 \o_buffer_reg[63][12]  (.D(n_123_76), .CK(n_120), .Q(
      \o_buffer[63] [12]), .QN());
   DFF_X1 \o_buffer_reg[63][11]  (.D(n_123_75), .CK(n_120), .Q(
      \o_buffer[63] [11]), .QN());
   DFF_X1 \o_buffer_reg[63][10]  (.D(n_123_74), .CK(n_120), .Q(
      \o_buffer[63] [10]), .QN());
   DFF_X1 \o_buffer_reg[63][9]  (.D(n_123_73), .CK(n_120), .Q(\o_buffer[63] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][8]  (.D(n_123_72), .CK(n_120), .Q(\o_buffer[63] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][7]  (.D(n_123_71), .CK(n_120), .Q(\o_buffer[63] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][6]  (.D(n_123_70), .CK(n_120), .Q(\o_buffer[63] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][5]  (.D(n_123_69), .CK(n_120), .Q(\o_buffer[63] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][4]  (.D(n_123_68), .CK(n_120), .Q(\o_buffer[63] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][3]  (.D(n_123_67), .CK(n_120), .Q(\o_buffer[63] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][2]  (.D(n_123_66), .CK(n_120), .Q(\o_buffer[63] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][1]  (.D(n_123_65), .CK(n_120), .Q(\o_buffer[63] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[63][0]  (.D(n_123_64), .CK(n_120), .Q(\o_buffer[63] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][15]  (.D(n_123_63), .CK(n_120), .Q(
      \o_buffer[62] [15]), .QN());
   DFF_X1 \o_buffer_reg[62][14]  (.D(n_123_62), .CK(n_120), .Q(
      \o_buffer[62] [14]), .QN());
   DFF_X1 \o_buffer_reg[62][13]  (.D(n_123_61), .CK(n_120), .Q(
      \o_buffer[62] [13]), .QN());
   DFF_X1 \o_buffer_reg[62][12]  (.D(n_123_60), .CK(n_120), .Q(
      \o_buffer[62] [12]), .QN());
   DFF_X1 \o_buffer_reg[62][11]  (.D(n_123_59), .CK(n_120), .Q(
      \o_buffer[62] [11]), .QN());
   DFF_X1 \o_buffer_reg[62][10]  (.D(n_123_58), .CK(n_120), .Q(
      \o_buffer[62] [10]), .QN());
   DFF_X1 \o_buffer_reg[62][9]  (.D(n_123_57), .CK(n_120), .Q(\o_buffer[62] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][8]  (.D(n_123_56), .CK(n_120), .Q(\o_buffer[62] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][7]  (.D(n_123_55), .CK(n_120), .Q(\o_buffer[62] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][6]  (.D(n_123_54), .CK(n_120), .Q(\o_buffer[62] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][5]  (.D(n_123_53), .CK(n_120), .Q(\o_buffer[62] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][4]  (.D(n_123_52), .CK(n_120), .Q(\o_buffer[62] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][3]  (.D(n_123_51), .CK(n_120), .Q(\o_buffer[62] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][2]  (.D(n_123_50), .CK(n_120), .Q(\o_buffer[62] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][1]  (.D(n_123_49), .CK(n_120), .Q(\o_buffer[62] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[62][0]  (.D(n_123_48), .CK(n_120), .Q(\o_buffer[62] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][15]  (.D(n_123_47), .CK(n_120), .Q(
      \o_buffer[61] [15]), .QN());
   DFF_X1 \o_buffer_reg[61][14]  (.D(n_123_46), .CK(n_120), .Q(
      \o_buffer[61] [14]), .QN());
   DFF_X1 \o_buffer_reg[61][13]  (.D(n_123_45), .CK(n_120), .Q(
      \o_buffer[61] [13]), .QN());
   DFF_X1 \o_buffer_reg[61][12]  (.D(n_123_44), .CK(n_120), .Q(
      \o_buffer[61] [12]), .QN());
   DFF_X1 \o_buffer_reg[61][11]  (.D(n_123_43), .CK(n_120), .Q(
      \o_buffer[61] [11]), .QN());
   DFF_X1 \o_buffer_reg[61][10]  (.D(n_123_42), .CK(n_120), .Q(
      \o_buffer[61] [10]), .QN());
   DFF_X1 \o_buffer_reg[61][9]  (.D(n_123_41), .CK(n_120), .Q(\o_buffer[61] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][8]  (.D(n_123_40), .CK(n_120), .Q(\o_buffer[61] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][7]  (.D(n_123_39), .CK(n_120), .Q(\o_buffer[61] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][6]  (.D(n_123_38), .CK(n_120), .Q(\o_buffer[61] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][5]  (.D(n_123_37), .CK(n_120), .Q(\o_buffer[61] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][4]  (.D(n_123_36), .CK(n_120), .Q(\o_buffer[61] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][3]  (.D(n_123_35), .CK(n_120), .Q(\o_buffer[61] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][2]  (.D(n_123_34), .CK(n_120), .Q(\o_buffer[61] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][1]  (.D(n_123_33), .CK(n_120), .Q(\o_buffer[61] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[61][0]  (.D(n_123_32), .CK(n_120), .Q(\o_buffer[61] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][15]  (.D(n_123_31), .CK(n_120), .Q(
      \o_buffer[60] [15]), .QN());
   DFF_X1 \o_buffer_reg[60][14]  (.D(n_123_30), .CK(n_120), .Q(
      \o_buffer[60] [14]), .QN());
   DFF_X1 \o_buffer_reg[60][13]  (.D(n_123_29), .CK(n_120), .Q(
      \o_buffer[60] [13]), .QN());
   DFF_X1 \o_buffer_reg[60][12]  (.D(n_123_28), .CK(n_120), .Q(
      \o_buffer[60] [12]), .QN());
   DFF_X1 \o_buffer_reg[60][11]  (.D(n_123_27), .CK(n_120), .Q(
      \o_buffer[60] [11]), .QN());
   DFF_X1 \o_buffer_reg[60][10]  (.D(n_123_26), .CK(n_120), .Q(
      \o_buffer[60] [10]), .QN());
   DFF_X1 \o_buffer_reg[60][9]  (.D(n_123_25), .CK(n_120), .Q(\o_buffer[60] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][8]  (.D(n_123_24), .CK(n_120), .Q(\o_buffer[60] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][7]  (.D(n_123_23), .CK(n_120), .Q(\o_buffer[60] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][6]  (.D(n_123_22), .CK(n_120), .Q(\o_buffer[60] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][5]  (.D(n_123_21), .CK(n_120), .Q(\o_buffer[60] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][4]  (.D(n_123_20), .CK(n_120), .Q(\o_buffer[60] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][3]  (.D(n_123_19), .CK(n_120), .Q(\o_buffer[60] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][2]  (.D(n_123_18), .CK(n_120), .Q(\o_buffer[60] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][1]  (.D(n_123_17), .CK(n_120), .Q(\o_buffer[60] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[60][0]  (.D(n_123_16), .CK(n_120), .Q(\o_buffer[60] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][15]  (.D(n_123_15), .CK(n_120), .Q(
      \o_buffer[59] [15]), .QN());
   DFF_X1 \o_buffer_reg[59][14]  (.D(n_123_14), .CK(n_120), .Q(
      \o_buffer[59] [14]), .QN());
   DFF_X1 \o_buffer_reg[59][13]  (.D(n_123_13), .CK(n_120), .Q(
      \o_buffer[59] [13]), .QN());
   DFF_X1 \o_buffer_reg[59][12]  (.D(n_123_12), .CK(n_120), .Q(
      \o_buffer[59] [12]), .QN());
   DFF_X1 \o_buffer_reg[59][11]  (.D(n_123_11), .CK(n_120), .Q(
      \o_buffer[59] [11]), .QN());
   DFF_X1 \o_buffer_reg[59][10]  (.D(n_123_10), .CK(n_120), .Q(
      \o_buffer[59] [10]), .QN());
   DFF_X1 \o_buffer_reg[59][9]  (.D(n_123_9), .CK(n_120), .Q(\o_buffer[59] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][8]  (.D(n_123_8), .CK(n_120), .Q(\o_buffer[59] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][7]  (.D(n_123_7), .CK(n_120), .Q(\o_buffer[59] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][6]  (.D(n_123_6), .CK(n_120), .Q(\o_buffer[59] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][5]  (.D(n_123_5), .CK(n_120), .Q(\o_buffer[59] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][4]  (.D(n_123_4), .CK(n_120), .Q(\o_buffer[59] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][3]  (.D(n_123_3), .CK(n_120), .Q(\o_buffer[59] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][2]  (.D(n_123_2), .CK(n_120), .Q(\o_buffer[59] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][1]  (.D(n_123_1), .CK(n_120), .Q(\o_buffer[59] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[59][0]  (.D(n_123_0), .CK(n_120), .Q(\o_buffer[59] [0]), 
      .QN());
   MUX2_X1 i_123_0_0 (.A(\o_buffer[118] [15]), .B(i_mem_data[15]), .S(n_1), 
      .Z(n_123_959));
   MUX2_X1 i_123_0_1 (.A(\o_buffer[118] [14]), .B(i_mem_data[14]), .S(n_1), 
      .Z(n_123_958));
   MUX2_X1 i_123_0_2 (.A(\o_buffer[118] [13]), .B(i_mem_data[13]), .S(n_1), 
      .Z(n_123_957));
   MUX2_X1 i_123_0_3 (.A(\o_buffer[118] [12]), .B(i_mem_data[12]), .S(n_1), 
      .Z(n_123_956));
   MUX2_X1 i_123_0_4 (.A(\o_buffer[118] [11]), .B(i_mem_data[11]), .S(n_1), 
      .Z(n_123_955));
   MUX2_X1 i_123_0_5 (.A(\o_buffer[118] [10]), .B(i_mem_data[10]), .S(n_1), 
      .Z(n_123_954));
   MUX2_X1 i_123_0_6 (.A(\o_buffer[118] [9]), .B(i_mem_data[9]), .S(n_1), 
      .Z(n_123_953));
   MUX2_X1 i_123_0_7 (.A(\o_buffer[118] [8]), .B(i_mem_data[8]), .S(n_1), 
      .Z(n_123_952));
   MUX2_X1 i_123_0_8 (.A(\o_buffer[118] [7]), .B(i_mem_data[7]), .S(n_1), 
      .Z(n_123_951));
   MUX2_X1 i_123_0_9 (.A(\o_buffer[118] [6]), .B(i_mem_data[6]), .S(n_1), 
      .Z(n_123_950));
   MUX2_X1 i_123_0_10 (.A(\o_buffer[118] [5]), .B(i_mem_data[5]), .S(n_1), 
      .Z(n_123_949));
   MUX2_X1 i_123_0_11 (.A(\o_buffer[118] [4]), .B(i_mem_data[4]), .S(n_1), 
      .Z(n_123_948));
   MUX2_X1 i_123_0_12 (.A(\o_buffer[118] [3]), .B(i_mem_data[3]), .S(n_1), 
      .Z(n_123_947));
   MUX2_X1 i_123_0_13 (.A(\o_buffer[118] [2]), .B(i_mem_data[2]), .S(n_1), 
      .Z(n_123_946));
   MUX2_X1 i_123_0_14 (.A(\o_buffer[118] [1]), .B(i_mem_data[1]), .S(n_1), 
      .Z(n_123_945));
   MUX2_X1 i_123_0_15 (.A(\o_buffer[118] [0]), .B(i_mem_data[0]), .S(n_1), 
      .Z(n_123_944));
   MUX2_X1 i_123_0_16 (.A(\o_buffer[117] [15]), .B(i_mem_data[15]), .S(n_2), 
      .Z(n_123_943));
   MUX2_X1 i_123_0_17 (.A(\o_buffer[117] [14]), .B(i_mem_data[14]), .S(n_2), 
      .Z(n_123_942));
   MUX2_X1 i_123_0_18 (.A(\o_buffer[117] [13]), .B(i_mem_data[13]), .S(n_2), 
      .Z(n_123_941));
   MUX2_X1 i_123_0_19 (.A(\o_buffer[117] [12]), .B(i_mem_data[12]), .S(n_2), 
      .Z(n_123_940));
   MUX2_X1 i_123_0_20 (.A(\o_buffer[117] [11]), .B(i_mem_data[11]), .S(n_2), 
      .Z(n_123_939));
   MUX2_X1 i_123_0_21 (.A(\o_buffer[117] [10]), .B(i_mem_data[10]), .S(n_2), 
      .Z(n_123_938));
   MUX2_X1 i_123_0_22 (.A(\o_buffer[117] [9]), .B(i_mem_data[9]), .S(n_2), 
      .Z(n_123_937));
   MUX2_X1 i_123_0_23 (.A(\o_buffer[117] [8]), .B(i_mem_data[8]), .S(n_2), 
      .Z(n_123_936));
   MUX2_X1 i_123_0_24 (.A(\o_buffer[117] [7]), .B(i_mem_data[7]), .S(n_2), 
      .Z(n_123_935));
   MUX2_X1 i_123_0_25 (.A(\o_buffer[117] [6]), .B(i_mem_data[6]), .S(n_2), 
      .Z(n_123_934));
   MUX2_X1 i_123_0_26 (.A(\o_buffer[117] [5]), .B(i_mem_data[5]), .S(n_2), 
      .Z(n_123_933));
   MUX2_X1 i_123_0_27 (.A(\o_buffer[117] [4]), .B(i_mem_data[4]), .S(n_2), 
      .Z(n_123_932));
   MUX2_X1 i_123_0_28 (.A(\o_buffer[117] [3]), .B(i_mem_data[3]), .S(n_2), 
      .Z(n_123_931));
   MUX2_X1 i_123_0_29 (.A(\o_buffer[117] [2]), .B(i_mem_data[2]), .S(n_2), 
      .Z(n_123_930));
   MUX2_X1 i_123_0_30 (.A(\o_buffer[117] [1]), .B(i_mem_data[1]), .S(n_2), 
      .Z(n_123_929));
   MUX2_X1 i_123_0_31 (.A(\o_buffer[117] [0]), .B(i_mem_data[0]), .S(n_2), 
      .Z(n_123_928));
   MUX2_X1 i_123_0_32 (.A(\o_buffer[116] [15]), .B(i_mem_data[15]), .S(n_3), 
      .Z(n_123_927));
   MUX2_X1 i_123_0_33 (.A(\o_buffer[116] [14]), .B(i_mem_data[14]), .S(n_3), 
      .Z(n_123_926));
   MUX2_X1 i_123_0_34 (.A(\o_buffer[116] [13]), .B(i_mem_data[13]), .S(n_3), 
      .Z(n_123_925));
   MUX2_X1 i_123_0_35 (.A(\o_buffer[116] [12]), .B(i_mem_data[12]), .S(n_3), 
      .Z(n_123_924));
   MUX2_X1 i_123_0_36 (.A(\o_buffer[116] [11]), .B(i_mem_data[11]), .S(n_3), 
      .Z(n_123_923));
   MUX2_X1 i_123_0_37 (.A(\o_buffer[116] [10]), .B(i_mem_data[10]), .S(n_3), 
      .Z(n_123_922));
   MUX2_X1 i_123_0_38 (.A(\o_buffer[116] [9]), .B(i_mem_data[9]), .S(n_3), 
      .Z(n_123_921));
   MUX2_X1 i_123_0_39 (.A(\o_buffer[116] [8]), .B(i_mem_data[8]), .S(n_3), 
      .Z(n_123_920));
   MUX2_X1 i_123_0_40 (.A(\o_buffer[116] [7]), .B(i_mem_data[7]), .S(n_3), 
      .Z(n_123_919));
   MUX2_X1 i_123_0_41 (.A(\o_buffer[116] [6]), .B(i_mem_data[6]), .S(n_3), 
      .Z(n_123_918));
   MUX2_X1 i_123_0_42 (.A(\o_buffer[116] [5]), .B(i_mem_data[5]), .S(n_3), 
      .Z(n_123_917));
   MUX2_X1 i_123_0_43 (.A(\o_buffer[116] [4]), .B(i_mem_data[4]), .S(n_3), 
      .Z(n_123_916));
   MUX2_X1 i_123_0_44 (.A(\o_buffer[116] [3]), .B(i_mem_data[3]), .S(n_3), 
      .Z(n_123_915));
   MUX2_X1 i_123_0_45 (.A(\o_buffer[116] [2]), .B(i_mem_data[2]), .S(n_3), 
      .Z(n_123_914));
   MUX2_X1 i_123_0_46 (.A(\o_buffer[116] [1]), .B(i_mem_data[1]), .S(n_3), 
      .Z(n_123_913));
   MUX2_X1 i_123_0_47 (.A(\o_buffer[116] [0]), .B(i_mem_data[0]), .S(n_3), 
      .Z(n_123_912));
   MUX2_X1 i_123_0_48 (.A(\o_buffer[115] [15]), .B(i_mem_data[15]), .S(n_4), 
      .Z(n_123_911));
   MUX2_X1 i_123_0_49 (.A(\o_buffer[115] [14]), .B(i_mem_data[14]), .S(n_4), 
      .Z(n_123_910));
   MUX2_X1 i_123_0_50 (.A(\o_buffer[115] [13]), .B(i_mem_data[13]), .S(n_4), 
      .Z(n_123_909));
   MUX2_X1 i_123_0_51 (.A(\o_buffer[115] [12]), .B(i_mem_data[12]), .S(n_4), 
      .Z(n_123_908));
   MUX2_X1 i_123_0_52 (.A(\o_buffer[115] [11]), .B(i_mem_data[11]), .S(n_4), 
      .Z(n_123_907));
   MUX2_X1 i_123_0_53 (.A(\o_buffer[115] [10]), .B(i_mem_data[10]), .S(n_4), 
      .Z(n_123_906));
   MUX2_X1 i_123_0_54 (.A(\o_buffer[115] [9]), .B(i_mem_data[9]), .S(n_4), 
      .Z(n_123_905));
   MUX2_X1 i_123_0_55 (.A(\o_buffer[115] [8]), .B(i_mem_data[8]), .S(n_4), 
      .Z(n_123_904));
   MUX2_X1 i_123_0_56 (.A(\o_buffer[115] [7]), .B(i_mem_data[7]), .S(n_4), 
      .Z(n_123_903));
   MUX2_X1 i_123_0_57 (.A(\o_buffer[115] [6]), .B(i_mem_data[6]), .S(n_4), 
      .Z(n_123_902));
   MUX2_X1 i_123_0_58 (.A(\o_buffer[115] [5]), .B(i_mem_data[5]), .S(n_4), 
      .Z(n_123_901));
   MUX2_X1 i_123_0_59 (.A(\o_buffer[115] [4]), .B(i_mem_data[4]), .S(n_4), 
      .Z(n_123_900));
   MUX2_X1 i_123_0_60 (.A(\o_buffer[115] [3]), .B(i_mem_data[3]), .S(n_4), 
      .Z(n_123_899));
   MUX2_X1 i_123_0_61 (.A(\o_buffer[115] [2]), .B(i_mem_data[2]), .S(n_4), 
      .Z(n_123_898));
   MUX2_X1 i_123_0_62 (.A(\o_buffer[115] [1]), .B(i_mem_data[1]), .S(n_4), 
      .Z(n_123_897));
   MUX2_X1 i_123_0_63 (.A(\o_buffer[115] [0]), .B(i_mem_data[0]), .S(n_4), 
      .Z(n_123_896));
   MUX2_X1 i_123_0_64 (.A(\o_buffer[114] [15]), .B(i_mem_data[15]), .S(n_5), 
      .Z(n_123_895));
   MUX2_X1 i_123_0_65 (.A(\o_buffer[114] [14]), .B(i_mem_data[14]), .S(n_5), 
      .Z(n_123_894));
   MUX2_X1 i_123_0_66 (.A(\o_buffer[114] [13]), .B(i_mem_data[13]), .S(n_5), 
      .Z(n_123_893));
   MUX2_X1 i_123_0_67 (.A(\o_buffer[114] [12]), .B(i_mem_data[12]), .S(n_5), 
      .Z(n_123_892));
   MUX2_X1 i_123_0_68 (.A(\o_buffer[114] [11]), .B(i_mem_data[11]), .S(n_5), 
      .Z(n_123_891));
   MUX2_X1 i_123_0_69 (.A(\o_buffer[114] [10]), .B(i_mem_data[10]), .S(n_5), 
      .Z(n_123_890));
   MUX2_X1 i_123_0_70 (.A(\o_buffer[114] [9]), .B(i_mem_data[9]), .S(n_5), 
      .Z(n_123_889));
   MUX2_X1 i_123_0_71 (.A(\o_buffer[114] [8]), .B(i_mem_data[8]), .S(n_5), 
      .Z(n_123_888));
   MUX2_X1 i_123_0_72 (.A(\o_buffer[114] [7]), .B(i_mem_data[7]), .S(n_5), 
      .Z(n_123_887));
   MUX2_X1 i_123_0_73 (.A(\o_buffer[114] [6]), .B(i_mem_data[6]), .S(n_5), 
      .Z(n_123_886));
   MUX2_X1 i_123_0_74 (.A(\o_buffer[114] [5]), .B(i_mem_data[5]), .S(n_5), 
      .Z(n_123_885));
   MUX2_X1 i_123_0_75 (.A(\o_buffer[114] [4]), .B(i_mem_data[4]), .S(n_5), 
      .Z(n_123_884));
   MUX2_X1 i_123_0_76 (.A(\o_buffer[114] [3]), .B(i_mem_data[3]), .S(n_5), 
      .Z(n_123_883));
   MUX2_X1 i_123_0_77 (.A(\o_buffer[114] [2]), .B(i_mem_data[2]), .S(n_5), 
      .Z(n_123_882));
   MUX2_X1 i_123_0_78 (.A(\o_buffer[114] [1]), .B(i_mem_data[1]), .S(n_5), 
      .Z(n_123_881));
   MUX2_X1 i_123_0_79 (.A(\o_buffer[114] [0]), .B(i_mem_data[0]), .S(n_5), 
      .Z(n_123_880));
   MUX2_X1 i_123_0_80 (.A(\o_buffer[113] [15]), .B(i_mem_data[15]), .S(n_6), 
      .Z(n_123_879));
   MUX2_X1 i_123_0_81 (.A(\o_buffer[113] [14]), .B(i_mem_data[14]), .S(n_6), 
      .Z(n_123_878));
   MUX2_X1 i_123_0_82 (.A(\o_buffer[113] [13]), .B(i_mem_data[13]), .S(n_6), 
      .Z(n_123_877));
   MUX2_X1 i_123_0_83 (.A(\o_buffer[113] [12]), .B(i_mem_data[12]), .S(n_6), 
      .Z(n_123_876));
   MUX2_X1 i_123_0_84 (.A(\o_buffer[113] [11]), .B(i_mem_data[11]), .S(n_6), 
      .Z(n_123_875));
   MUX2_X1 i_123_0_85 (.A(\o_buffer[113] [10]), .B(i_mem_data[10]), .S(n_6), 
      .Z(n_123_874));
   MUX2_X1 i_123_0_86 (.A(\o_buffer[113] [9]), .B(i_mem_data[9]), .S(n_6), 
      .Z(n_123_873));
   MUX2_X1 i_123_0_87 (.A(\o_buffer[113] [8]), .B(i_mem_data[8]), .S(n_6), 
      .Z(n_123_872));
   MUX2_X1 i_123_0_88 (.A(\o_buffer[113] [7]), .B(i_mem_data[7]), .S(n_6), 
      .Z(n_123_871));
   MUX2_X1 i_123_0_89 (.A(\o_buffer[113] [6]), .B(i_mem_data[6]), .S(n_6), 
      .Z(n_123_870));
   MUX2_X1 i_123_0_90 (.A(\o_buffer[113] [5]), .B(i_mem_data[5]), .S(n_6), 
      .Z(n_123_869));
   MUX2_X1 i_123_0_91 (.A(\o_buffer[113] [4]), .B(i_mem_data[4]), .S(n_6), 
      .Z(n_123_868));
   MUX2_X1 i_123_0_92 (.A(\o_buffer[113] [3]), .B(i_mem_data[3]), .S(n_6), 
      .Z(n_123_867));
   MUX2_X1 i_123_0_93 (.A(\o_buffer[113] [2]), .B(i_mem_data[2]), .S(n_6), 
      .Z(n_123_866));
   MUX2_X1 i_123_0_94 (.A(\o_buffer[113] [1]), .B(i_mem_data[1]), .S(n_6), 
      .Z(n_123_865));
   MUX2_X1 i_123_0_95 (.A(\o_buffer[113] [0]), .B(i_mem_data[0]), .S(n_6), 
      .Z(n_123_864));
   MUX2_X1 i_123_0_96 (.A(\o_buffer[112] [15]), .B(i_mem_data[15]), .S(n_7), 
      .Z(n_123_863));
   MUX2_X1 i_123_0_97 (.A(\o_buffer[112] [14]), .B(i_mem_data[14]), .S(n_7), 
      .Z(n_123_862));
   MUX2_X1 i_123_0_98 (.A(\o_buffer[112] [13]), .B(i_mem_data[13]), .S(n_7), 
      .Z(n_123_861));
   MUX2_X1 i_123_0_99 (.A(\o_buffer[112] [12]), .B(i_mem_data[12]), .S(n_7), 
      .Z(n_123_860));
   MUX2_X1 i_123_0_100 (.A(\o_buffer[112] [11]), .B(i_mem_data[11]), .S(n_7), 
      .Z(n_123_859));
   MUX2_X1 i_123_0_101 (.A(\o_buffer[112] [10]), .B(i_mem_data[10]), .S(n_7), 
      .Z(n_123_858));
   MUX2_X1 i_123_0_102 (.A(\o_buffer[112] [9]), .B(i_mem_data[9]), .S(n_7), 
      .Z(n_123_857));
   MUX2_X1 i_123_0_103 (.A(\o_buffer[112] [8]), .B(i_mem_data[8]), .S(n_7), 
      .Z(n_123_856));
   MUX2_X1 i_123_0_104 (.A(\o_buffer[112] [7]), .B(i_mem_data[7]), .S(n_7), 
      .Z(n_123_855));
   MUX2_X1 i_123_0_105 (.A(\o_buffer[112] [6]), .B(i_mem_data[6]), .S(n_7), 
      .Z(n_123_854));
   MUX2_X1 i_123_0_106 (.A(\o_buffer[112] [5]), .B(i_mem_data[5]), .S(n_7), 
      .Z(n_123_853));
   MUX2_X1 i_123_0_107 (.A(\o_buffer[112] [4]), .B(i_mem_data[4]), .S(n_7), 
      .Z(n_123_852));
   MUX2_X1 i_123_0_108 (.A(\o_buffer[112] [3]), .B(i_mem_data[3]), .S(n_7), 
      .Z(n_123_851));
   MUX2_X1 i_123_0_109 (.A(\o_buffer[112] [2]), .B(i_mem_data[2]), .S(n_7), 
      .Z(n_123_850));
   MUX2_X1 i_123_0_110 (.A(\o_buffer[112] [1]), .B(i_mem_data[1]), .S(n_7), 
      .Z(n_123_849));
   MUX2_X1 i_123_0_111 (.A(\o_buffer[112] [0]), .B(i_mem_data[0]), .S(n_7), 
      .Z(n_123_848));
   MUX2_X1 i_123_0_112 (.A(\o_buffer[111] [15]), .B(i_mem_data[15]), .S(n_8), 
      .Z(n_123_847));
   MUX2_X1 i_123_0_113 (.A(\o_buffer[111] [14]), .B(i_mem_data[14]), .S(n_8), 
      .Z(n_123_846));
   MUX2_X1 i_123_0_114 (.A(\o_buffer[111] [13]), .B(i_mem_data[13]), .S(n_8), 
      .Z(n_123_845));
   MUX2_X1 i_123_0_115 (.A(\o_buffer[111] [12]), .B(i_mem_data[12]), .S(n_8), 
      .Z(n_123_844));
   MUX2_X1 i_123_0_116 (.A(\o_buffer[111] [11]), .B(i_mem_data[11]), .S(n_8), 
      .Z(n_123_843));
   MUX2_X1 i_123_0_117 (.A(\o_buffer[111] [10]), .B(i_mem_data[10]), .S(n_8), 
      .Z(n_123_842));
   MUX2_X1 i_123_0_118 (.A(\o_buffer[111] [9]), .B(i_mem_data[9]), .S(n_8), 
      .Z(n_123_841));
   MUX2_X1 i_123_0_119 (.A(\o_buffer[111] [8]), .B(i_mem_data[8]), .S(n_8), 
      .Z(n_123_840));
   MUX2_X1 i_123_0_120 (.A(\o_buffer[111] [7]), .B(i_mem_data[7]), .S(n_8), 
      .Z(n_123_839));
   MUX2_X1 i_123_0_121 (.A(\o_buffer[111] [6]), .B(i_mem_data[6]), .S(n_8), 
      .Z(n_123_838));
   MUX2_X1 i_123_0_122 (.A(\o_buffer[111] [5]), .B(i_mem_data[5]), .S(n_8), 
      .Z(n_123_837));
   MUX2_X1 i_123_0_123 (.A(\o_buffer[111] [4]), .B(i_mem_data[4]), .S(n_8), 
      .Z(n_123_836));
   MUX2_X1 i_123_0_124 (.A(\o_buffer[111] [3]), .B(i_mem_data[3]), .S(n_8), 
      .Z(n_123_835));
   MUX2_X1 i_123_0_125 (.A(\o_buffer[111] [2]), .B(i_mem_data[2]), .S(n_8), 
      .Z(n_123_834));
   MUX2_X1 i_123_0_126 (.A(\o_buffer[111] [1]), .B(i_mem_data[1]), .S(n_8), 
      .Z(n_123_833));
   MUX2_X1 i_123_0_127 (.A(\o_buffer[111] [0]), .B(i_mem_data[0]), .S(n_8), 
      .Z(n_123_832));
   MUX2_X1 i_123_0_128 (.A(\o_buffer[110] [15]), .B(i_mem_data[15]), .S(n_9), 
      .Z(n_123_831));
   MUX2_X1 i_123_0_129 (.A(\o_buffer[110] [14]), .B(i_mem_data[14]), .S(n_9), 
      .Z(n_123_830));
   MUX2_X1 i_123_0_130 (.A(\o_buffer[110] [13]), .B(i_mem_data[13]), .S(n_9), 
      .Z(n_123_829));
   MUX2_X1 i_123_0_131 (.A(\o_buffer[110] [12]), .B(i_mem_data[12]), .S(n_9), 
      .Z(n_123_828));
   MUX2_X1 i_123_0_132 (.A(\o_buffer[110] [11]), .B(i_mem_data[11]), .S(n_9), 
      .Z(n_123_827));
   MUX2_X1 i_123_0_133 (.A(\o_buffer[110] [10]), .B(i_mem_data[10]), .S(n_9), 
      .Z(n_123_826));
   MUX2_X1 i_123_0_134 (.A(\o_buffer[110] [9]), .B(i_mem_data[9]), .S(n_9), 
      .Z(n_123_825));
   MUX2_X1 i_123_0_135 (.A(\o_buffer[110] [8]), .B(i_mem_data[8]), .S(n_9), 
      .Z(n_123_824));
   MUX2_X1 i_123_0_136 (.A(\o_buffer[110] [7]), .B(i_mem_data[7]), .S(n_9), 
      .Z(n_123_823));
   MUX2_X1 i_123_0_137 (.A(\o_buffer[110] [6]), .B(i_mem_data[6]), .S(n_9), 
      .Z(n_123_822));
   MUX2_X1 i_123_0_138 (.A(\o_buffer[110] [5]), .B(i_mem_data[5]), .S(n_9), 
      .Z(n_123_821));
   MUX2_X1 i_123_0_139 (.A(\o_buffer[110] [4]), .B(i_mem_data[4]), .S(n_9), 
      .Z(n_123_820));
   MUX2_X1 i_123_0_140 (.A(\o_buffer[110] [3]), .B(i_mem_data[3]), .S(n_9), 
      .Z(n_123_819));
   MUX2_X1 i_123_0_141 (.A(\o_buffer[110] [2]), .B(i_mem_data[2]), .S(n_9), 
      .Z(n_123_818));
   MUX2_X1 i_123_0_142 (.A(\o_buffer[110] [1]), .B(i_mem_data[1]), .S(n_9), 
      .Z(n_123_817));
   MUX2_X1 i_123_0_143 (.A(\o_buffer[110] [0]), .B(i_mem_data[0]), .S(n_9), 
      .Z(n_123_816));
   MUX2_X1 i_123_0_144 (.A(\o_buffer[109] [15]), .B(i_mem_data[15]), .S(n_10), 
      .Z(n_123_815));
   MUX2_X1 i_123_0_145 (.A(\o_buffer[109] [14]), .B(i_mem_data[14]), .S(n_10), 
      .Z(n_123_814));
   MUX2_X1 i_123_0_146 (.A(\o_buffer[109] [13]), .B(i_mem_data[13]), .S(n_10), 
      .Z(n_123_813));
   MUX2_X1 i_123_0_147 (.A(\o_buffer[109] [12]), .B(i_mem_data[12]), .S(n_10), 
      .Z(n_123_812));
   MUX2_X1 i_123_0_148 (.A(\o_buffer[109] [11]), .B(i_mem_data[11]), .S(n_10), 
      .Z(n_123_811));
   MUX2_X1 i_123_0_149 (.A(\o_buffer[109] [10]), .B(i_mem_data[10]), .S(n_10), 
      .Z(n_123_810));
   MUX2_X1 i_123_0_150 (.A(\o_buffer[109] [9]), .B(i_mem_data[9]), .S(n_10), 
      .Z(n_123_809));
   MUX2_X1 i_123_0_151 (.A(\o_buffer[109] [8]), .B(i_mem_data[8]), .S(n_10), 
      .Z(n_123_808));
   MUX2_X1 i_123_0_152 (.A(\o_buffer[109] [7]), .B(i_mem_data[7]), .S(n_10), 
      .Z(n_123_807));
   MUX2_X1 i_123_0_153 (.A(\o_buffer[109] [6]), .B(i_mem_data[6]), .S(n_10), 
      .Z(n_123_806));
   MUX2_X1 i_123_0_154 (.A(\o_buffer[109] [5]), .B(i_mem_data[5]), .S(n_10), 
      .Z(n_123_805));
   MUX2_X1 i_123_0_155 (.A(\o_buffer[109] [4]), .B(i_mem_data[4]), .S(n_10), 
      .Z(n_123_804));
   MUX2_X1 i_123_0_156 (.A(\o_buffer[109] [3]), .B(i_mem_data[3]), .S(n_10), 
      .Z(n_123_803));
   MUX2_X1 i_123_0_157 (.A(\o_buffer[109] [2]), .B(i_mem_data[2]), .S(n_10), 
      .Z(n_123_802));
   MUX2_X1 i_123_0_158 (.A(\o_buffer[109] [1]), .B(i_mem_data[1]), .S(n_10), 
      .Z(n_123_801));
   MUX2_X1 i_123_0_159 (.A(\o_buffer[109] [0]), .B(i_mem_data[0]), .S(n_10), 
      .Z(n_123_800));
   MUX2_X1 i_123_0_160 (.A(\o_buffer[108] [15]), .B(i_mem_data[15]), .S(n_11), 
      .Z(n_123_799));
   MUX2_X1 i_123_0_161 (.A(\o_buffer[108] [14]), .B(i_mem_data[14]), .S(n_11), 
      .Z(n_123_798));
   MUX2_X1 i_123_0_162 (.A(\o_buffer[108] [13]), .B(i_mem_data[13]), .S(n_11), 
      .Z(n_123_797));
   MUX2_X1 i_123_0_163 (.A(\o_buffer[108] [12]), .B(i_mem_data[12]), .S(n_11), 
      .Z(n_123_796));
   MUX2_X1 i_123_0_164 (.A(\o_buffer[108] [11]), .B(i_mem_data[11]), .S(n_11), 
      .Z(n_123_795));
   MUX2_X1 i_123_0_165 (.A(\o_buffer[108] [10]), .B(i_mem_data[10]), .S(n_11), 
      .Z(n_123_794));
   MUX2_X1 i_123_0_166 (.A(\o_buffer[108] [9]), .B(i_mem_data[9]), .S(n_11), 
      .Z(n_123_793));
   MUX2_X1 i_123_0_167 (.A(\o_buffer[108] [8]), .B(i_mem_data[8]), .S(n_11), 
      .Z(n_123_792));
   MUX2_X1 i_123_0_168 (.A(\o_buffer[108] [7]), .B(i_mem_data[7]), .S(n_11), 
      .Z(n_123_791));
   MUX2_X1 i_123_0_169 (.A(\o_buffer[108] [6]), .B(i_mem_data[6]), .S(n_11), 
      .Z(n_123_790));
   MUX2_X1 i_123_0_170 (.A(\o_buffer[108] [5]), .B(i_mem_data[5]), .S(n_11), 
      .Z(n_123_789));
   MUX2_X1 i_123_0_171 (.A(\o_buffer[108] [4]), .B(i_mem_data[4]), .S(n_11), 
      .Z(n_123_788));
   MUX2_X1 i_123_0_172 (.A(\o_buffer[108] [3]), .B(i_mem_data[3]), .S(n_11), 
      .Z(n_123_787));
   MUX2_X1 i_123_0_173 (.A(\o_buffer[108] [2]), .B(i_mem_data[2]), .S(n_11), 
      .Z(n_123_786));
   MUX2_X1 i_123_0_174 (.A(\o_buffer[108] [1]), .B(i_mem_data[1]), .S(n_11), 
      .Z(n_123_785));
   MUX2_X1 i_123_0_175 (.A(\o_buffer[108] [0]), .B(i_mem_data[0]), .S(n_11), 
      .Z(n_123_784));
   MUX2_X1 i_123_0_176 (.A(\o_buffer[107] [15]), .B(i_mem_data[15]), .S(n_12), 
      .Z(n_123_783));
   MUX2_X1 i_123_0_177 (.A(\o_buffer[107] [14]), .B(i_mem_data[14]), .S(n_12), 
      .Z(n_123_782));
   MUX2_X1 i_123_0_178 (.A(\o_buffer[107] [13]), .B(i_mem_data[13]), .S(n_12), 
      .Z(n_123_781));
   MUX2_X1 i_123_0_179 (.A(\o_buffer[107] [12]), .B(i_mem_data[12]), .S(n_12), 
      .Z(n_123_780));
   MUX2_X1 i_123_0_180 (.A(\o_buffer[107] [11]), .B(i_mem_data[11]), .S(n_12), 
      .Z(n_123_779));
   MUX2_X1 i_123_0_181 (.A(\o_buffer[107] [10]), .B(i_mem_data[10]), .S(n_12), 
      .Z(n_123_778));
   MUX2_X1 i_123_0_182 (.A(\o_buffer[107] [9]), .B(i_mem_data[9]), .S(n_12), 
      .Z(n_123_777));
   MUX2_X1 i_123_0_183 (.A(\o_buffer[107] [8]), .B(i_mem_data[8]), .S(n_12), 
      .Z(n_123_776));
   MUX2_X1 i_123_0_184 (.A(\o_buffer[107] [7]), .B(i_mem_data[7]), .S(n_12), 
      .Z(n_123_775));
   MUX2_X1 i_123_0_185 (.A(\o_buffer[107] [6]), .B(i_mem_data[6]), .S(n_12), 
      .Z(n_123_774));
   MUX2_X1 i_123_0_186 (.A(\o_buffer[107] [5]), .B(i_mem_data[5]), .S(n_12), 
      .Z(n_123_773));
   MUX2_X1 i_123_0_187 (.A(\o_buffer[107] [4]), .B(i_mem_data[4]), .S(n_12), 
      .Z(n_123_772));
   MUX2_X1 i_123_0_188 (.A(\o_buffer[107] [3]), .B(i_mem_data[3]), .S(n_12), 
      .Z(n_123_771));
   MUX2_X1 i_123_0_189 (.A(\o_buffer[107] [2]), .B(i_mem_data[2]), .S(n_12), 
      .Z(n_123_770));
   MUX2_X1 i_123_0_190 (.A(\o_buffer[107] [1]), .B(i_mem_data[1]), .S(n_12), 
      .Z(n_123_769));
   MUX2_X1 i_123_0_191 (.A(\o_buffer[107] [0]), .B(i_mem_data[0]), .S(n_12), 
      .Z(n_123_768));
   MUX2_X1 i_123_0_192 (.A(\o_buffer[106] [15]), .B(i_mem_data[15]), .S(n_13), 
      .Z(n_123_767));
   MUX2_X1 i_123_0_193 (.A(\o_buffer[106] [14]), .B(i_mem_data[14]), .S(n_13), 
      .Z(n_123_766));
   MUX2_X1 i_123_0_194 (.A(\o_buffer[106] [13]), .B(i_mem_data[13]), .S(n_13), 
      .Z(n_123_765));
   MUX2_X1 i_123_0_195 (.A(\o_buffer[106] [12]), .B(i_mem_data[12]), .S(n_13), 
      .Z(n_123_764));
   MUX2_X1 i_123_0_196 (.A(\o_buffer[106] [11]), .B(i_mem_data[11]), .S(n_13), 
      .Z(n_123_763));
   MUX2_X1 i_123_0_197 (.A(\o_buffer[106] [10]), .B(i_mem_data[10]), .S(n_13), 
      .Z(n_123_762));
   MUX2_X1 i_123_0_198 (.A(\o_buffer[106] [9]), .B(i_mem_data[9]), .S(n_13), 
      .Z(n_123_761));
   MUX2_X1 i_123_0_199 (.A(\o_buffer[106] [8]), .B(i_mem_data[8]), .S(n_13), 
      .Z(n_123_760));
   MUX2_X1 i_123_0_200 (.A(\o_buffer[106] [7]), .B(i_mem_data[7]), .S(n_13), 
      .Z(n_123_759));
   MUX2_X1 i_123_0_201 (.A(\o_buffer[106] [6]), .B(i_mem_data[6]), .S(n_13), 
      .Z(n_123_758));
   MUX2_X1 i_123_0_202 (.A(\o_buffer[106] [5]), .B(i_mem_data[5]), .S(n_13), 
      .Z(n_123_757));
   MUX2_X1 i_123_0_203 (.A(\o_buffer[106] [4]), .B(i_mem_data[4]), .S(n_13), 
      .Z(n_123_756));
   MUX2_X1 i_123_0_204 (.A(\o_buffer[106] [3]), .B(i_mem_data[3]), .S(n_13), 
      .Z(n_123_755));
   MUX2_X1 i_123_0_205 (.A(\o_buffer[106] [2]), .B(i_mem_data[2]), .S(n_13), 
      .Z(n_123_754));
   MUX2_X1 i_123_0_206 (.A(\o_buffer[106] [1]), .B(i_mem_data[1]), .S(n_13), 
      .Z(n_123_753));
   MUX2_X1 i_123_0_207 (.A(\o_buffer[106] [0]), .B(i_mem_data[0]), .S(n_13), 
      .Z(n_123_752));
   MUX2_X1 i_123_0_208 (.A(\o_buffer[105] [15]), .B(i_mem_data[15]), .S(n_14), 
      .Z(n_123_751));
   MUX2_X1 i_123_0_209 (.A(\o_buffer[105] [14]), .B(i_mem_data[14]), .S(n_14), 
      .Z(n_123_750));
   MUX2_X1 i_123_0_210 (.A(\o_buffer[105] [13]), .B(i_mem_data[13]), .S(n_14), 
      .Z(n_123_749));
   MUX2_X1 i_123_0_211 (.A(\o_buffer[105] [12]), .B(i_mem_data[12]), .S(n_14), 
      .Z(n_123_748));
   MUX2_X1 i_123_0_212 (.A(\o_buffer[105] [11]), .B(i_mem_data[11]), .S(n_14), 
      .Z(n_123_747));
   MUX2_X1 i_123_0_213 (.A(\o_buffer[105] [10]), .B(i_mem_data[10]), .S(n_14), 
      .Z(n_123_746));
   MUX2_X1 i_123_0_214 (.A(\o_buffer[105] [9]), .B(i_mem_data[9]), .S(n_14), 
      .Z(n_123_745));
   MUX2_X1 i_123_0_215 (.A(\o_buffer[105] [8]), .B(i_mem_data[8]), .S(n_14), 
      .Z(n_123_744));
   MUX2_X1 i_123_0_216 (.A(\o_buffer[105] [7]), .B(i_mem_data[7]), .S(n_14), 
      .Z(n_123_743));
   MUX2_X1 i_123_0_217 (.A(\o_buffer[105] [6]), .B(i_mem_data[6]), .S(n_14), 
      .Z(n_123_742));
   MUX2_X1 i_123_0_218 (.A(\o_buffer[105] [5]), .B(i_mem_data[5]), .S(n_14), 
      .Z(n_123_741));
   MUX2_X1 i_123_0_219 (.A(\o_buffer[105] [4]), .B(i_mem_data[4]), .S(n_14), 
      .Z(n_123_740));
   MUX2_X1 i_123_0_220 (.A(\o_buffer[105] [3]), .B(i_mem_data[3]), .S(n_14), 
      .Z(n_123_739));
   MUX2_X1 i_123_0_221 (.A(\o_buffer[105] [2]), .B(i_mem_data[2]), .S(n_14), 
      .Z(n_123_738));
   MUX2_X1 i_123_0_222 (.A(\o_buffer[105] [1]), .B(i_mem_data[1]), .S(n_14), 
      .Z(n_123_737));
   MUX2_X1 i_123_0_223 (.A(\o_buffer[105] [0]), .B(i_mem_data[0]), .S(n_14), 
      .Z(n_123_736));
   MUX2_X1 i_123_0_224 (.A(\o_buffer[104] [15]), .B(i_mem_data[15]), .S(n_15), 
      .Z(n_123_735));
   MUX2_X1 i_123_0_225 (.A(\o_buffer[104] [14]), .B(i_mem_data[14]), .S(n_15), 
      .Z(n_123_734));
   MUX2_X1 i_123_0_226 (.A(\o_buffer[104] [13]), .B(i_mem_data[13]), .S(n_15), 
      .Z(n_123_733));
   MUX2_X1 i_123_0_227 (.A(\o_buffer[104] [12]), .B(i_mem_data[12]), .S(n_15), 
      .Z(n_123_732));
   MUX2_X1 i_123_0_228 (.A(\o_buffer[104] [11]), .B(i_mem_data[11]), .S(n_15), 
      .Z(n_123_731));
   MUX2_X1 i_123_0_229 (.A(\o_buffer[104] [10]), .B(i_mem_data[10]), .S(n_15), 
      .Z(n_123_730));
   MUX2_X1 i_123_0_230 (.A(\o_buffer[104] [9]), .B(i_mem_data[9]), .S(n_15), 
      .Z(n_123_729));
   MUX2_X1 i_123_0_231 (.A(\o_buffer[104] [8]), .B(i_mem_data[8]), .S(n_15), 
      .Z(n_123_728));
   MUX2_X1 i_123_0_232 (.A(\o_buffer[104] [7]), .B(i_mem_data[7]), .S(n_15), 
      .Z(n_123_727));
   MUX2_X1 i_123_0_233 (.A(\o_buffer[104] [6]), .B(i_mem_data[6]), .S(n_15), 
      .Z(n_123_726));
   MUX2_X1 i_123_0_234 (.A(\o_buffer[104] [5]), .B(i_mem_data[5]), .S(n_15), 
      .Z(n_123_725));
   MUX2_X1 i_123_0_235 (.A(\o_buffer[104] [4]), .B(i_mem_data[4]), .S(n_15), 
      .Z(n_123_724));
   MUX2_X1 i_123_0_236 (.A(\o_buffer[104] [3]), .B(i_mem_data[3]), .S(n_15), 
      .Z(n_123_723));
   MUX2_X1 i_123_0_237 (.A(\o_buffer[104] [2]), .B(i_mem_data[2]), .S(n_15), 
      .Z(n_123_722));
   MUX2_X1 i_123_0_238 (.A(\o_buffer[104] [1]), .B(i_mem_data[1]), .S(n_15), 
      .Z(n_123_721));
   MUX2_X1 i_123_0_239 (.A(\o_buffer[104] [0]), .B(i_mem_data[0]), .S(n_15), 
      .Z(n_123_720));
   MUX2_X1 i_123_0_240 (.A(\o_buffer[103] [15]), .B(i_mem_data[15]), .S(n_16), 
      .Z(n_123_719));
   MUX2_X1 i_123_0_241 (.A(\o_buffer[103] [14]), .B(i_mem_data[14]), .S(n_16), 
      .Z(n_123_718));
   MUX2_X1 i_123_0_242 (.A(\o_buffer[103] [13]), .B(i_mem_data[13]), .S(n_16), 
      .Z(n_123_717));
   MUX2_X1 i_123_0_243 (.A(\o_buffer[103] [12]), .B(i_mem_data[12]), .S(n_16), 
      .Z(n_123_716));
   MUX2_X1 i_123_0_244 (.A(\o_buffer[103] [11]), .B(i_mem_data[11]), .S(n_16), 
      .Z(n_123_715));
   MUX2_X1 i_123_0_245 (.A(\o_buffer[103] [10]), .B(i_mem_data[10]), .S(n_16), 
      .Z(n_123_714));
   MUX2_X1 i_123_0_246 (.A(\o_buffer[103] [9]), .B(i_mem_data[9]), .S(n_16), 
      .Z(n_123_713));
   MUX2_X1 i_123_0_247 (.A(\o_buffer[103] [8]), .B(i_mem_data[8]), .S(n_16), 
      .Z(n_123_712));
   MUX2_X1 i_123_0_248 (.A(\o_buffer[103] [7]), .B(i_mem_data[7]), .S(n_16), 
      .Z(n_123_711));
   MUX2_X1 i_123_0_249 (.A(\o_buffer[103] [6]), .B(i_mem_data[6]), .S(n_16), 
      .Z(n_123_710));
   MUX2_X1 i_123_0_250 (.A(\o_buffer[103] [5]), .B(i_mem_data[5]), .S(n_16), 
      .Z(n_123_709));
   MUX2_X1 i_123_0_251 (.A(\o_buffer[103] [4]), .B(i_mem_data[4]), .S(n_16), 
      .Z(n_123_708));
   MUX2_X1 i_123_0_252 (.A(\o_buffer[103] [3]), .B(i_mem_data[3]), .S(n_16), 
      .Z(n_123_707));
   MUX2_X1 i_123_0_253 (.A(\o_buffer[103] [2]), .B(i_mem_data[2]), .S(n_16), 
      .Z(n_123_706));
   MUX2_X1 i_123_0_254 (.A(\o_buffer[103] [1]), .B(i_mem_data[1]), .S(n_16), 
      .Z(n_123_705));
   MUX2_X1 i_123_0_255 (.A(\o_buffer[103] [0]), .B(i_mem_data[0]), .S(n_16), 
      .Z(n_123_704));
   MUX2_X1 i_123_0_256 (.A(\o_buffer[102] [15]), .B(i_mem_data[15]), .S(n_17), 
      .Z(n_123_703));
   MUX2_X1 i_123_0_257 (.A(\o_buffer[102] [14]), .B(i_mem_data[14]), .S(n_17), 
      .Z(n_123_702));
   MUX2_X1 i_123_0_258 (.A(\o_buffer[102] [13]), .B(i_mem_data[13]), .S(n_17), 
      .Z(n_123_701));
   MUX2_X1 i_123_0_259 (.A(\o_buffer[102] [12]), .B(i_mem_data[12]), .S(n_17), 
      .Z(n_123_700));
   MUX2_X1 i_123_0_260 (.A(\o_buffer[102] [11]), .B(i_mem_data[11]), .S(n_17), 
      .Z(n_123_699));
   MUX2_X1 i_123_0_261 (.A(\o_buffer[102] [10]), .B(i_mem_data[10]), .S(n_17), 
      .Z(n_123_698));
   MUX2_X1 i_123_0_262 (.A(\o_buffer[102] [9]), .B(i_mem_data[9]), .S(n_17), 
      .Z(n_123_697));
   MUX2_X1 i_123_0_263 (.A(\o_buffer[102] [8]), .B(i_mem_data[8]), .S(n_17), 
      .Z(n_123_696));
   MUX2_X1 i_123_0_264 (.A(\o_buffer[102] [7]), .B(i_mem_data[7]), .S(n_17), 
      .Z(n_123_695));
   MUX2_X1 i_123_0_265 (.A(\o_buffer[102] [6]), .B(i_mem_data[6]), .S(n_17), 
      .Z(n_123_694));
   MUX2_X1 i_123_0_266 (.A(\o_buffer[102] [5]), .B(i_mem_data[5]), .S(n_17), 
      .Z(n_123_693));
   MUX2_X1 i_123_0_267 (.A(\o_buffer[102] [4]), .B(i_mem_data[4]), .S(n_17), 
      .Z(n_123_692));
   MUX2_X1 i_123_0_268 (.A(\o_buffer[102] [3]), .B(i_mem_data[3]), .S(n_17), 
      .Z(n_123_691));
   MUX2_X1 i_123_0_269 (.A(\o_buffer[102] [2]), .B(i_mem_data[2]), .S(n_17), 
      .Z(n_123_690));
   MUX2_X1 i_123_0_270 (.A(\o_buffer[102] [1]), .B(i_mem_data[1]), .S(n_17), 
      .Z(n_123_689));
   MUX2_X1 i_123_0_271 (.A(\o_buffer[102] [0]), .B(i_mem_data[0]), .S(n_17), 
      .Z(n_123_688));
   MUX2_X1 i_123_0_272 (.A(\o_buffer[101] [15]), .B(i_mem_data[15]), .S(n_18), 
      .Z(n_123_687));
   MUX2_X1 i_123_0_273 (.A(\o_buffer[101] [14]), .B(i_mem_data[14]), .S(n_18), 
      .Z(n_123_686));
   MUX2_X1 i_123_0_274 (.A(\o_buffer[101] [13]), .B(i_mem_data[13]), .S(n_18), 
      .Z(n_123_685));
   MUX2_X1 i_123_0_275 (.A(\o_buffer[101] [12]), .B(i_mem_data[12]), .S(n_18), 
      .Z(n_123_684));
   MUX2_X1 i_123_0_276 (.A(\o_buffer[101] [11]), .B(i_mem_data[11]), .S(n_18), 
      .Z(n_123_683));
   MUX2_X1 i_123_0_277 (.A(\o_buffer[101] [10]), .B(i_mem_data[10]), .S(n_18), 
      .Z(n_123_682));
   MUX2_X1 i_123_0_278 (.A(\o_buffer[101] [9]), .B(i_mem_data[9]), .S(n_18), 
      .Z(n_123_681));
   MUX2_X1 i_123_0_279 (.A(\o_buffer[101] [8]), .B(i_mem_data[8]), .S(n_18), 
      .Z(n_123_680));
   MUX2_X1 i_123_0_280 (.A(\o_buffer[101] [7]), .B(i_mem_data[7]), .S(n_18), 
      .Z(n_123_679));
   MUX2_X1 i_123_0_281 (.A(\o_buffer[101] [6]), .B(i_mem_data[6]), .S(n_18), 
      .Z(n_123_678));
   MUX2_X1 i_123_0_282 (.A(\o_buffer[101] [5]), .B(i_mem_data[5]), .S(n_18), 
      .Z(n_123_677));
   MUX2_X1 i_123_0_283 (.A(\o_buffer[101] [4]), .B(i_mem_data[4]), .S(n_18), 
      .Z(n_123_676));
   MUX2_X1 i_123_0_284 (.A(\o_buffer[101] [3]), .B(i_mem_data[3]), .S(n_18), 
      .Z(n_123_675));
   MUX2_X1 i_123_0_285 (.A(\o_buffer[101] [2]), .B(i_mem_data[2]), .S(n_18), 
      .Z(n_123_674));
   MUX2_X1 i_123_0_286 (.A(\o_buffer[101] [1]), .B(i_mem_data[1]), .S(n_18), 
      .Z(n_123_673));
   MUX2_X1 i_123_0_287 (.A(\o_buffer[101] [0]), .B(i_mem_data[0]), .S(n_18), 
      .Z(n_123_672));
   MUX2_X1 i_123_0_288 (.A(\o_buffer[100] [15]), .B(i_mem_data[15]), .S(n_19), 
      .Z(n_123_671));
   MUX2_X1 i_123_0_289 (.A(\o_buffer[100] [14]), .B(i_mem_data[14]), .S(n_19), 
      .Z(n_123_670));
   MUX2_X1 i_123_0_290 (.A(\o_buffer[100] [13]), .B(i_mem_data[13]), .S(n_19), 
      .Z(n_123_669));
   MUX2_X1 i_123_0_291 (.A(\o_buffer[100] [12]), .B(i_mem_data[12]), .S(n_19), 
      .Z(n_123_668));
   MUX2_X1 i_123_0_292 (.A(\o_buffer[100] [11]), .B(i_mem_data[11]), .S(n_19), 
      .Z(n_123_667));
   MUX2_X1 i_123_0_293 (.A(\o_buffer[100] [10]), .B(i_mem_data[10]), .S(n_19), 
      .Z(n_123_666));
   MUX2_X1 i_123_0_294 (.A(\o_buffer[100] [9]), .B(i_mem_data[9]), .S(n_19), 
      .Z(n_123_665));
   MUX2_X1 i_123_0_295 (.A(\o_buffer[100] [8]), .B(i_mem_data[8]), .S(n_19), 
      .Z(n_123_664));
   MUX2_X1 i_123_0_296 (.A(\o_buffer[100] [7]), .B(i_mem_data[7]), .S(n_19), 
      .Z(n_123_663));
   MUX2_X1 i_123_0_297 (.A(\o_buffer[100] [6]), .B(i_mem_data[6]), .S(n_19), 
      .Z(n_123_662));
   MUX2_X1 i_123_0_298 (.A(\o_buffer[100] [5]), .B(i_mem_data[5]), .S(n_19), 
      .Z(n_123_661));
   MUX2_X1 i_123_0_299 (.A(\o_buffer[100] [4]), .B(i_mem_data[4]), .S(n_19), 
      .Z(n_123_660));
   MUX2_X1 i_123_0_300 (.A(\o_buffer[100] [3]), .B(i_mem_data[3]), .S(n_19), 
      .Z(n_123_659));
   MUX2_X1 i_123_0_301 (.A(\o_buffer[100] [2]), .B(i_mem_data[2]), .S(n_19), 
      .Z(n_123_658));
   MUX2_X1 i_123_0_302 (.A(\o_buffer[100] [1]), .B(i_mem_data[1]), .S(n_19), 
      .Z(n_123_657));
   MUX2_X1 i_123_0_303 (.A(\o_buffer[100] [0]), .B(i_mem_data[0]), .S(n_19), 
      .Z(n_123_656));
   MUX2_X1 i_123_0_304 (.A(\o_buffer[99] [15]), .B(i_mem_data[15]), .S(n_20), 
      .Z(n_123_655));
   MUX2_X1 i_123_0_305 (.A(\o_buffer[99] [14]), .B(i_mem_data[14]), .S(n_20), 
      .Z(n_123_654));
   MUX2_X1 i_123_0_306 (.A(\o_buffer[99] [13]), .B(i_mem_data[13]), .S(n_20), 
      .Z(n_123_653));
   MUX2_X1 i_123_0_307 (.A(\o_buffer[99] [12]), .B(i_mem_data[12]), .S(n_20), 
      .Z(n_123_652));
   MUX2_X1 i_123_0_308 (.A(\o_buffer[99] [11]), .B(i_mem_data[11]), .S(n_20), 
      .Z(n_123_651));
   MUX2_X1 i_123_0_309 (.A(\o_buffer[99] [10]), .B(i_mem_data[10]), .S(n_20), 
      .Z(n_123_650));
   MUX2_X1 i_123_0_310 (.A(\o_buffer[99] [9]), .B(i_mem_data[9]), .S(n_20), 
      .Z(n_123_649));
   MUX2_X1 i_123_0_311 (.A(\o_buffer[99] [8]), .B(i_mem_data[8]), .S(n_20), 
      .Z(n_123_648));
   MUX2_X1 i_123_0_312 (.A(\o_buffer[99] [7]), .B(i_mem_data[7]), .S(n_20), 
      .Z(n_123_647));
   MUX2_X1 i_123_0_313 (.A(\o_buffer[99] [6]), .B(i_mem_data[6]), .S(n_20), 
      .Z(n_123_646));
   MUX2_X1 i_123_0_314 (.A(\o_buffer[99] [5]), .B(i_mem_data[5]), .S(n_20), 
      .Z(n_123_645));
   MUX2_X1 i_123_0_315 (.A(\o_buffer[99] [4]), .B(i_mem_data[4]), .S(n_20), 
      .Z(n_123_644));
   MUX2_X1 i_123_0_316 (.A(\o_buffer[99] [3]), .B(i_mem_data[3]), .S(n_20), 
      .Z(n_123_643));
   MUX2_X1 i_123_0_317 (.A(\o_buffer[99] [2]), .B(i_mem_data[2]), .S(n_20), 
      .Z(n_123_642));
   MUX2_X1 i_123_0_318 (.A(\o_buffer[99] [1]), .B(i_mem_data[1]), .S(n_20), 
      .Z(n_123_641));
   MUX2_X1 i_123_0_319 (.A(\o_buffer[99] [0]), .B(i_mem_data[0]), .S(n_20), 
      .Z(n_123_640));
   MUX2_X1 i_123_0_320 (.A(\o_buffer[98] [15]), .B(i_mem_data[15]), .S(n_21), 
      .Z(n_123_639));
   MUX2_X1 i_123_0_321 (.A(\o_buffer[98] [14]), .B(i_mem_data[14]), .S(n_21), 
      .Z(n_123_638));
   MUX2_X1 i_123_0_322 (.A(\o_buffer[98] [13]), .B(i_mem_data[13]), .S(n_21), 
      .Z(n_123_637));
   MUX2_X1 i_123_0_323 (.A(\o_buffer[98] [12]), .B(i_mem_data[12]), .S(n_21), 
      .Z(n_123_636));
   MUX2_X1 i_123_0_324 (.A(\o_buffer[98] [11]), .B(i_mem_data[11]), .S(n_21), 
      .Z(n_123_635));
   MUX2_X1 i_123_0_325 (.A(\o_buffer[98] [10]), .B(i_mem_data[10]), .S(n_21), 
      .Z(n_123_634));
   MUX2_X1 i_123_0_326 (.A(\o_buffer[98] [9]), .B(i_mem_data[9]), .S(n_21), 
      .Z(n_123_633));
   MUX2_X1 i_123_0_327 (.A(\o_buffer[98] [8]), .B(i_mem_data[8]), .S(n_21), 
      .Z(n_123_632));
   MUX2_X1 i_123_0_328 (.A(\o_buffer[98] [7]), .B(i_mem_data[7]), .S(n_21), 
      .Z(n_123_631));
   MUX2_X1 i_123_0_329 (.A(\o_buffer[98] [6]), .B(i_mem_data[6]), .S(n_21), 
      .Z(n_123_630));
   MUX2_X1 i_123_0_330 (.A(\o_buffer[98] [5]), .B(i_mem_data[5]), .S(n_21), 
      .Z(n_123_629));
   MUX2_X1 i_123_0_331 (.A(\o_buffer[98] [4]), .B(i_mem_data[4]), .S(n_21), 
      .Z(n_123_628));
   MUX2_X1 i_123_0_332 (.A(\o_buffer[98] [3]), .B(i_mem_data[3]), .S(n_21), 
      .Z(n_123_627));
   MUX2_X1 i_123_0_333 (.A(\o_buffer[98] [2]), .B(i_mem_data[2]), .S(n_21), 
      .Z(n_123_626));
   MUX2_X1 i_123_0_334 (.A(\o_buffer[98] [1]), .B(i_mem_data[1]), .S(n_21), 
      .Z(n_123_625));
   MUX2_X1 i_123_0_335 (.A(\o_buffer[98] [0]), .B(i_mem_data[0]), .S(n_21), 
      .Z(n_123_624));
   MUX2_X1 i_123_0_336 (.A(\o_buffer[97] [15]), .B(i_mem_data[15]), .S(n_22), 
      .Z(n_123_623));
   MUX2_X1 i_123_0_337 (.A(\o_buffer[97] [14]), .B(i_mem_data[14]), .S(n_22), 
      .Z(n_123_622));
   MUX2_X1 i_123_0_338 (.A(\o_buffer[97] [13]), .B(i_mem_data[13]), .S(n_22), 
      .Z(n_123_621));
   MUX2_X1 i_123_0_339 (.A(\o_buffer[97] [12]), .B(i_mem_data[12]), .S(n_22), 
      .Z(n_123_620));
   MUX2_X1 i_123_0_340 (.A(\o_buffer[97] [11]), .B(i_mem_data[11]), .S(n_22), 
      .Z(n_123_619));
   MUX2_X1 i_123_0_341 (.A(\o_buffer[97] [10]), .B(i_mem_data[10]), .S(n_22), 
      .Z(n_123_618));
   MUX2_X1 i_123_0_342 (.A(\o_buffer[97] [9]), .B(i_mem_data[9]), .S(n_22), 
      .Z(n_123_617));
   MUX2_X1 i_123_0_343 (.A(\o_buffer[97] [8]), .B(i_mem_data[8]), .S(n_22), 
      .Z(n_123_616));
   MUX2_X1 i_123_0_344 (.A(\o_buffer[97] [7]), .B(i_mem_data[7]), .S(n_22), 
      .Z(n_123_615));
   MUX2_X1 i_123_0_345 (.A(\o_buffer[97] [6]), .B(i_mem_data[6]), .S(n_22), 
      .Z(n_123_614));
   MUX2_X1 i_123_0_346 (.A(\o_buffer[97] [5]), .B(i_mem_data[5]), .S(n_22), 
      .Z(n_123_613));
   MUX2_X1 i_123_0_347 (.A(\o_buffer[97] [4]), .B(i_mem_data[4]), .S(n_22), 
      .Z(n_123_612));
   MUX2_X1 i_123_0_348 (.A(\o_buffer[97] [3]), .B(i_mem_data[3]), .S(n_22), 
      .Z(n_123_611));
   MUX2_X1 i_123_0_349 (.A(\o_buffer[97] [2]), .B(i_mem_data[2]), .S(n_22), 
      .Z(n_123_610));
   MUX2_X1 i_123_0_350 (.A(\o_buffer[97] [1]), .B(i_mem_data[1]), .S(n_22), 
      .Z(n_123_609));
   MUX2_X1 i_123_0_351 (.A(\o_buffer[97] [0]), .B(i_mem_data[0]), .S(n_22), 
      .Z(n_123_608));
   MUX2_X1 i_123_0_352 (.A(\o_buffer[96] [15]), .B(i_mem_data[15]), .S(n_23), 
      .Z(n_123_607));
   MUX2_X1 i_123_0_353 (.A(\o_buffer[96] [14]), .B(i_mem_data[14]), .S(n_23), 
      .Z(n_123_606));
   MUX2_X1 i_123_0_354 (.A(\o_buffer[96] [13]), .B(i_mem_data[13]), .S(n_23), 
      .Z(n_123_605));
   MUX2_X1 i_123_0_355 (.A(\o_buffer[96] [12]), .B(i_mem_data[12]), .S(n_23), 
      .Z(n_123_604));
   MUX2_X1 i_123_0_356 (.A(\o_buffer[96] [11]), .B(i_mem_data[11]), .S(n_23), 
      .Z(n_123_603));
   MUX2_X1 i_123_0_357 (.A(\o_buffer[96] [10]), .B(i_mem_data[10]), .S(n_23), 
      .Z(n_123_602));
   MUX2_X1 i_123_0_358 (.A(\o_buffer[96] [9]), .B(i_mem_data[9]), .S(n_23), 
      .Z(n_123_601));
   MUX2_X1 i_123_0_359 (.A(\o_buffer[96] [8]), .B(i_mem_data[8]), .S(n_23), 
      .Z(n_123_600));
   MUX2_X1 i_123_0_360 (.A(\o_buffer[96] [7]), .B(i_mem_data[7]), .S(n_23), 
      .Z(n_123_599));
   MUX2_X1 i_123_0_361 (.A(\o_buffer[96] [6]), .B(i_mem_data[6]), .S(n_23), 
      .Z(n_123_598));
   MUX2_X1 i_123_0_362 (.A(\o_buffer[96] [5]), .B(i_mem_data[5]), .S(n_23), 
      .Z(n_123_597));
   MUX2_X1 i_123_0_363 (.A(\o_buffer[96] [4]), .B(i_mem_data[4]), .S(n_23), 
      .Z(n_123_596));
   MUX2_X1 i_123_0_364 (.A(\o_buffer[96] [3]), .B(i_mem_data[3]), .S(n_23), 
      .Z(n_123_595));
   MUX2_X1 i_123_0_365 (.A(\o_buffer[96] [2]), .B(i_mem_data[2]), .S(n_23), 
      .Z(n_123_594));
   MUX2_X1 i_123_0_366 (.A(\o_buffer[96] [1]), .B(i_mem_data[1]), .S(n_23), 
      .Z(n_123_593));
   MUX2_X1 i_123_0_367 (.A(\o_buffer[96] [0]), .B(i_mem_data[0]), .S(n_23), 
      .Z(n_123_592));
   MUX2_X1 i_123_0_368 (.A(\o_buffer[95] [15]), .B(i_mem_data[15]), .S(n_24), 
      .Z(n_123_591));
   MUX2_X1 i_123_0_369 (.A(\o_buffer[95] [14]), .B(i_mem_data[14]), .S(n_24), 
      .Z(n_123_590));
   MUX2_X1 i_123_0_370 (.A(\o_buffer[95] [13]), .B(i_mem_data[13]), .S(n_24), 
      .Z(n_123_589));
   MUX2_X1 i_123_0_371 (.A(\o_buffer[95] [12]), .B(i_mem_data[12]), .S(n_24), 
      .Z(n_123_588));
   MUX2_X1 i_123_0_372 (.A(\o_buffer[95] [11]), .B(i_mem_data[11]), .S(n_24), 
      .Z(n_123_587));
   MUX2_X1 i_123_0_373 (.A(\o_buffer[95] [10]), .B(i_mem_data[10]), .S(n_24), 
      .Z(n_123_586));
   MUX2_X1 i_123_0_374 (.A(\o_buffer[95] [9]), .B(i_mem_data[9]), .S(n_24), 
      .Z(n_123_585));
   MUX2_X1 i_123_0_375 (.A(\o_buffer[95] [8]), .B(i_mem_data[8]), .S(n_24), 
      .Z(n_123_584));
   MUX2_X1 i_123_0_376 (.A(\o_buffer[95] [7]), .B(i_mem_data[7]), .S(n_24), 
      .Z(n_123_583));
   MUX2_X1 i_123_0_377 (.A(\o_buffer[95] [6]), .B(i_mem_data[6]), .S(n_24), 
      .Z(n_123_582));
   MUX2_X1 i_123_0_378 (.A(\o_buffer[95] [5]), .B(i_mem_data[5]), .S(n_24), 
      .Z(n_123_581));
   MUX2_X1 i_123_0_379 (.A(\o_buffer[95] [4]), .B(i_mem_data[4]), .S(n_24), 
      .Z(n_123_580));
   MUX2_X1 i_123_0_380 (.A(\o_buffer[95] [3]), .B(i_mem_data[3]), .S(n_24), 
      .Z(n_123_579));
   MUX2_X1 i_123_0_381 (.A(\o_buffer[95] [2]), .B(i_mem_data[2]), .S(n_24), 
      .Z(n_123_578));
   MUX2_X1 i_123_0_382 (.A(\o_buffer[95] [1]), .B(i_mem_data[1]), .S(n_24), 
      .Z(n_123_577));
   MUX2_X1 i_123_0_383 (.A(\o_buffer[95] [0]), .B(i_mem_data[0]), .S(n_24), 
      .Z(n_123_576));
   MUX2_X1 i_123_0_384 (.A(\o_buffer[94] [15]), .B(i_mem_data[15]), .S(n_25), 
      .Z(n_123_575));
   MUX2_X1 i_123_0_385 (.A(\o_buffer[94] [14]), .B(i_mem_data[14]), .S(n_25), 
      .Z(n_123_574));
   MUX2_X1 i_123_0_386 (.A(\o_buffer[94] [13]), .B(i_mem_data[13]), .S(n_25), 
      .Z(n_123_573));
   MUX2_X1 i_123_0_387 (.A(\o_buffer[94] [12]), .B(i_mem_data[12]), .S(n_25), 
      .Z(n_123_572));
   MUX2_X1 i_123_0_388 (.A(\o_buffer[94] [11]), .B(i_mem_data[11]), .S(n_25), 
      .Z(n_123_571));
   MUX2_X1 i_123_0_389 (.A(\o_buffer[94] [10]), .B(i_mem_data[10]), .S(n_25), 
      .Z(n_123_570));
   MUX2_X1 i_123_0_390 (.A(\o_buffer[94] [9]), .B(i_mem_data[9]), .S(n_25), 
      .Z(n_123_569));
   MUX2_X1 i_123_0_391 (.A(\o_buffer[94] [8]), .B(i_mem_data[8]), .S(n_25), 
      .Z(n_123_568));
   MUX2_X1 i_123_0_392 (.A(\o_buffer[94] [7]), .B(i_mem_data[7]), .S(n_25), 
      .Z(n_123_567));
   MUX2_X1 i_123_0_393 (.A(\o_buffer[94] [6]), .B(i_mem_data[6]), .S(n_25), 
      .Z(n_123_566));
   MUX2_X1 i_123_0_394 (.A(\o_buffer[94] [5]), .B(i_mem_data[5]), .S(n_25), 
      .Z(n_123_565));
   MUX2_X1 i_123_0_395 (.A(\o_buffer[94] [4]), .B(i_mem_data[4]), .S(n_25), 
      .Z(n_123_564));
   MUX2_X1 i_123_0_396 (.A(\o_buffer[94] [3]), .B(i_mem_data[3]), .S(n_25), 
      .Z(n_123_563));
   MUX2_X1 i_123_0_397 (.A(\o_buffer[94] [2]), .B(i_mem_data[2]), .S(n_25), 
      .Z(n_123_562));
   MUX2_X1 i_123_0_398 (.A(\o_buffer[94] [1]), .B(i_mem_data[1]), .S(n_25), 
      .Z(n_123_561));
   MUX2_X1 i_123_0_399 (.A(\o_buffer[94] [0]), .B(i_mem_data[0]), .S(n_25), 
      .Z(n_123_560));
   MUX2_X1 i_123_0_400 (.A(\o_buffer[93] [15]), .B(i_mem_data[15]), .S(n_26), 
      .Z(n_123_559));
   MUX2_X1 i_123_0_401 (.A(\o_buffer[93] [14]), .B(i_mem_data[14]), .S(n_26), 
      .Z(n_123_558));
   MUX2_X1 i_123_0_402 (.A(\o_buffer[93] [13]), .B(i_mem_data[13]), .S(n_26), 
      .Z(n_123_557));
   MUX2_X1 i_123_0_403 (.A(\o_buffer[93] [12]), .B(i_mem_data[12]), .S(n_26), 
      .Z(n_123_556));
   MUX2_X1 i_123_0_404 (.A(\o_buffer[93] [11]), .B(i_mem_data[11]), .S(n_26), 
      .Z(n_123_555));
   MUX2_X1 i_123_0_405 (.A(\o_buffer[93] [10]), .B(i_mem_data[10]), .S(n_26), 
      .Z(n_123_554));
   MUX2_X1 i_123_0_406 (.A(\o_buffer[93] [9]), .B(i_mem_data[9]), .S(n_26), 
      .Z(n_123_553));
   MUX2_X1 i_123_0_407 (.A(\o_buffer[93] [8]), .B(i_mem_data[8]), .S(n_26), 
      .Z(n_123_552));
   MUX2_X1 i_123_0_408 (.A(\o_buffer[93] [7]), .B(i_mem_data[7]), .S(n_26), 
      .Z(n_123_551));
   MUX2_X1 i_123_0_409 (.A(\o_buffer[93] [6]), .B(i_mem_data[6]), .S(n_26), 
      .Z(n_123_550));
   MUX2_X1 i_123_0_410 (.A(\o_buffer[93] [5]), .B(i_mem_data[5]), .S(n_26), 
      .Z(n_123_549));
   MUX2_X1 i_123_0_411 (.A(\o_buffer[93] [4]), .B(i_mem_data[4]), .S(n_26), 
      .Z(n_123_548));
   MUX2_X1 i_123_0_412 (.A(\o_buffer[93] [3]), .B(i_mem_data[3]), .S(n_26), 
      .Z(n_123_547));
   MUX2_X1 i_123_0_413 (.A(\o_buffer[93] [2]), .B(i_mem_data[2]), .S(n_26), 
      .Z(n_123_546));
   MUX2_X1 i_123_0_414 (.A(\o_buffer[93] [1]), .B(i_mem_data[1]), .S(n_26), 
      .Z(n_123_545));
   MUX2_X1 i_123_0_415 (.A(\o_buffer[93] [0]), .B(i_mem_data[0]), .S(n_26), 
      .Z(n_123_544));
   MUX2_X1 i_123_0_416 (.A(\o_buffer[92] [15]), .B(i_mem_data[15]), .S(n_27), 
      .Z(n_123_543));
   MUX2_X1 i_123_0_417 (.A(\o_buffer[92] [14]), .B(i_mem_data[14]), .S(n_27), 
      .Z(n_123_542));
   MUX2_X1 i_123_0_418 (.A(\o_buffer[92] [13]), .B(i_mem_data[13]), .S(n_27), 
      .Z(n_123_541));
   MUX2_X1 i_123_0_419 (.A(\o_buffer[92] [12]), .B(i_mem_data[12]), .S(n_27), 
      .Z(n_123_540));
   MUX2_X1 i_123_0_420 (.A(\o_buffer[92] [11]), .B(i_mem_data[11]), .S(n_27), 
      .Z(n_123_539));
   MUX2_X1 i_123_0_421 (.A(\o_buffer[92] [10]), .B(i_mem_data[10]), .S(n_27), 
      .Z(n_123_538));
   MUX2_X1 i_123_0_422 (.A(\o_buffer[92] [9]), .B(i_mem_data[9]), .S(n_27), 
      .Z(n_123_537));
   MUX2_X1 i_123_0_423 (.A(\o_buffer[92] [8]), .B(i_mem_data[8]), .S(n_27), 
      .Z(n_123_536));
   MUX2_X1 i_123_0_424 (.A(\o_buffer[92] [7]), .B(i_mem_data[7]), .S(n_27), 
      .Z(n_123_535));
   MUX2_X1 i_123_0_425 (.A(\o_buffer[92] [6]), .B(i_mem_data[6]), .S(n_27), 
      .Z(n_123_534));
   MUX2_X1 i_123_0_426 (.A(\o_buffer[92] [5]), .B(i_mem_data[5]), .S(n_27), 
      .Z(n_123_533));
   MUX2_X1 i_123_0_427 (.A(\o_buffer[92] [4]), .B(i_mem_data[4]), .S(n_27), 
      .Z(n_123_532));
   MUX2_X1 i_123_0_428 (.A(\o_buffer[92] [3]), .B(i_mem_data[3]), .S(n_27), 
      .Z(n_123_531));
   MUX2_X1 i_123_0_429 (.A(\o_buffer[92] [2]), .B(i_mem_data[2]), .S(n_27), 
      .Z(n_123_530));
   MUX2_X1 i_123_0_430 (.A(\o_buffer[92] [1]), .B(i_mem_data[1]), .S(n_27), 
      .Z(n_123_529));
   MUX2_X1 i_123_0_431 (.A(\o_buffer[92] [0]), .B(i_mem_data[0]), .S(n_27), 
      .Z(n_123_528));
   MUX2_X1 i_123_0_432 (.A(\o_buffer[91] [15]), .B(i_mem_data[15]), .S(n_28), 
      .Z(n_123_527));
   MUX2_X1 i_123_0_433 (.A(\o_buffer[91] [14]), .B(i_mem_data[14]), .S(n_28), 
      .Z(n_123_526));
   MUX2_X1 i_123_0_434 (.A(\o_buffer[91] [13]), .B(i_mem_data[13]), .S(n_28), 
      .Z(n_123_525));
   MUX2_X1 i_123_0_435 (.A(\o_buffer[91] [12]), .B(i_mem_data[12]), .S(n_28), 
      .Z(n_123_524));
   MUX2_X1 i_123_0_436 (.A(\o_buffer[91] [11]), .B(i_mem_data[11]), .S(n_28), 
      .Z(n_123_523));
   MUX2_X1 i_123_0_437 (.A(\o_buffer[91] [10]), .B(i_mem_data[10]), .S(n_28), 
      .Z(n_123_522));
   MUX2_X1 i_123_0_438 (.A(\o_buffer[91] [9]), .B(i_mem_data[9]), .S(n_28), 
      .Z(n_123_521));
   MUX2_X1 i_123_0_439 (.A(\o_buffer[91] [8]), .B(i_mem_data[8]), .S(n_28), 
      .Z(n_123_520));
   MUX2_X1 i_123_0_440 (.A(\o_buffer[91] [7]), .B(i_mem_data[7]), .S(n_28), 
      .Z(n_123_519));
   MUX2_X1 i_123_0_441 (.A(\o_buffer[91] [6]), .B(i_mem_data[6]), .S(n_28), 
      .Z(n_123_518));
   MUX2_X1 i_123_0_442 (.A(\o_buffer[91] [5]), .B(i_mem_data[5]), .S(n_28), 
      .Z(n_123_517));
   MUX2_X1 i_123_0_443 (.A(\o_buffer[91] [4]), .B(i_mem_data[4]), .S(n_28), 
      .Z(n_123_516));
   MUX2_X1 i_123_0_444 (.A(\o_buffer[91] [3]), .B(i_mem_data[3]), .S(n_28), 
      .Z(n_123_515));
   MUX2_X1 i_123_0_445 (.A(\o_buffer[91] [2]), .B(i_mem_data[2]), .S(n_28), 
      .Z(n_123_514));
   MUX2_X1 i_123_0_446 (.A(\o_buffer[91] [1]), .B(i_mem_data[1]), .S(n_28), 
      .Z(n_123_513));
   MUX2_X1 i_123_0_447 (.A(\o_buffer[91] [0]), .B(i_mem_data[0]), .S(n_28), 
      .Z(n_123_512));
   MUX2_X1 i_123_0_448 (.A(\o_buffer[90] [15]), .B(i_mem_data[15]), .S(n_29), 
      .Z(n_123_511));
   MUX2_X1 i_123_0_449 (.A(\o_buffer[90] [14]), .B(i_mem_data[14]), .S(n_29), 
      .Z(n_123_510));
   MUX2_X1 i_123_0_450 (.A(\o_buffer[90] [13]), .B(i_mem_data[13]), .S(n_29), 
      .Z(n_123_509));
   MUX2_X1 i_123_0_451 (.A(\o_buffer[90] [12]), .B(i_mem_data[12]), .S(n_29), 
      .Z(n_123_508));
   MUX2_X1 i_123_0_452 (.A(\o_buffer[90] [11]), .B(i_mem_data[11]), .S(n_29), 
      .Z(n_123_507));
   MUX2_X1 i_123_0_453 (.A(\o_buffer[90] [10]), .B(i_mem_data[10]), .S(n_29), 
      .Z(n_123_506));
   MUX2_X1 i_123_0_454 (.A(\o_buffer[90] [9]), .B(i_mem_data[9]), .S(n_29), 
      .Z(n_123_505));
   MUX2_X1 i_123_0_455 (.A(\o_buffer[90] [8]), .B(i_mem_data[8]), .S(n_29), 
      .Z(n_123_504));
   MUX2_X1 i_123_0_456 (.A(\o_buffer[90] [7]), .B(i_mem_data[7]), .S(n_29), 
      .Z(n_123_503));
   MUX2_X1 i_123_0_457 (.A(\o_buffer[90] [6]), .B(i_mem_data[6]), .S(n_29), 
      .Z(n_123_502));
   MUX2_X1 i_123_0_458 (.A(\o_buffer[90] [5]), .B(i_mem_data[5]), .S(n_29), 
      .Z(n_123_501));
   MUX2_X1 i_123_0_459 (.A(\o_buffer[90] [4]), .B(i_mem_data[4]), .S(n_29), 
      .Z(n_123_500));
   MUX2_X1 i_123_0_460 (.A(\o_buffer[90] [3]), .B(i_mem_data[3]), .S(n_29), 
      .Z(n_123_499));
   MUX2_X1 i_123_0_461 (.A(\o_buffer[90] [2]), .B(i_mem_data[2]), .S(n_29), 
      .Z(n_123_498));
   MUX2_X1 i_123_0_462 (.A(\o_buffer[90] [1]), .B(i_mem_data[1]), .S(n_29), 
      .Z(n_123_497));
   MUX2_X1 i_123_0_463 (.A(\o_buffer[90] [0]), .B(i_mem_data[0]), .S(n_29), 
      .Z(n_123_496));
   MUX2_X1 i_123_0_464 (.A(\o_buffer[89] [15]), .B(i_mem_data[15]), .S(n_30), 
      .Z(n_123_495));
   MUX2_X1 i_123_0_465 (.A(\o_buffer[89] [14]), .B(i_mem_data[14]), .S(n_30), 
      .Z(n_123_494));
   MUX2_X1 i_123_0_466 (.A(\o_buffer[89] [13]), .B(i_mem_data[13]), .S(n_30), 
      .Z(n_123_493));
   MUX2_X1 i_123_0_467 (.A(\o_buffer[89] [12]), .B(i_mem_data[12]), .S(n_30), 
      .Z(n_123_492));
   MUX2_X1 i_123_0_468 (.A(\o_buffer[89] [11]), .B(i_mem_data[11]), .S(n_30), 
      .Z(n_123_491));
   MUX2_X1 i_123_0_469 (.A(\o_buffer[89] [10]), .B(i_mem_data[10]), .S(n_30), 
      .Z(n_123_490));
   MUX2_X1 i_123_0_470 (.A(\o_buffer[89] [9]), .B(i_mem_data[9]), .S(n_30), 
      .Z(n_123_489));
   MUX2_X1 i_123_0_471 (.A(\o_buffer[89] [8]), .B(i_mem_data[8]), .S(n_30), 
      .Z(n_123_488));
   MUX2_X1 i_123_0_472 (.A(\o_buffer[89] [7]), .B(i_mem_data[7]), .S(n_30), 
      .Z(n_123_487));
   MUX2_X1 i_123_0_473 (.A(\o_buffer[89] [6]), .B(i_mem_data[6]), .S(n_30), 
      .Z(n_123_486));
   MUX2_X1 i_123_0_474 (.A(\o_buffer[89] [5]), .B(i_mem_data[5]), .S(n_30), 
      .Z(n_123_485));
   MUX2_X1 i_123_0_475 (.A(\o_buffer[89] [4]), .B(i_mem_data[4]), .S(n_30), 
      .Z(n_123_484));
   MUX2_X1 i_123_0_476 (.A(\o_buffer[89] [3]), .B(i_mem_data[3]), .S(n_30), 
      .Z(n_123_483));
   MUX2_X1 i_123_0_477 (.A(\o_buffer[89] [2]), .B(i_mem_data[2]), .S(n_30), 
      .Z(n_123_482));
   MUX2_X1 i_123_0_478 (.A(\o_buffer[89] [1]), .B(i_mem_data[1]), .S(n_30), 
      .Z(n_123_481));
   MUX2_X1 i_123_0_479 (.A(\o_buffer[89] [0]), .B(i_mem_data[0]), .S(n_30), 
      .Z(n_123_480));
   MUX2_X1 i_123_0_480 (.A(\o_buffer[88] [15]), .B(i_mem_data[15]), .S(n_31), 
      .Z(n_123_479));
   MUX2_X1 i_123_0_481 (.A(\o_buffer[88] [14]), .B(i_mem_data[14]), .S(n_31), 
      .Z(n_123_478));
   MUX2_X1 i_123_0_482 (.A(\o_buffer[88] [13]), .B(i_mem_data[13]), .S(n_31), 
      .Z(n_123_477));
   MUX2_X1 i_123_0_483 (.A(\o_buffer[88] [12]), .B(i_mem_data[12]), .S(n_31), 
      .Z(n_123_476));
   MUX2_X1 i_123_0_484 (.A(\o_buffer[88] [11]), .B(i_mem_data[11]), .S(n_31), 
      .Z(n_123_475));
   MUX2_X1 i_123_0_485 (.A(\o_buffer[88] [10]), .B(i_mem_data[10]), .S(n_31), 
      .Z(n_123_474));
   MUX2_X1 i_123_0_486 (.A(\o_buffer[88] [9]), .B(i_mem_data[9]), .S(n_31), 
      .Z(n_123_473));
   MUX2_X1 i_123_0_487 (.A(\o_buffer[88] [8]), .B(i_mem_data[8]), .S(n_31), 
      .Z(n_123_472));
   MUX2_X1 i_123_0_488 (.A(\o_buffer[88] [7]), .B(i_mem_data[7]), .S(n_31), 
      .Z(n_123_471));
   MUX2_X1 i_123_0_489 (.A(\o_buffer[88] [6]), .B(i_mem_data[6]), .S(n_31), 
      .Z(n_123_470));
   MUX2_X1 i_123_0_490 (.A(\o_buffer[88] [5]), .B(i_mem_data[5]), .S(n_31), 
      .Z(n_123_469));
   MUX2_X1 i_123_0_491 (.A(\o_buffer[88] [4]), .B(i_mem_data[4]), .S(n_31), 
      .Z(n_123_468));
   MUX2_X1 i_123_0_492 (.A(\o_buffer[88] [3]), .B(i_mem_data[3]), .S(n_31), 
      .Z(n_123_467));
   MUX2_X1 i_123_0_493 (.A(\o_buffer[88] [2]), .B(i_mem_data[2]), .S(n_31), 
      .Z(n_123_466));
   MUX2_X1 i_123_0_494 (.A(\o_buffer[88] [1]), .B(i_mem_data[1]), .S(n_31), 
      .Z(n_123_465));
   MUX2_X1 i_123_0_495 (.A(\o_buffer[88] [0]), .B(i_mem_data[0]), .S(n_31), 
      .Z(n_123_464));
   MUX2_X1 i_123_0_496 (.A(\o_buffer[87] [15]), .B(i_mem_data[15]), .S(n_32), 
      .Z(n_123_463));
   MUX2_X1 i_123_0_497 (.A(\o_buffer[87] [14]), .B(i_mem_data[14]), .S(n_32), 
      .Z(n_123_462));
   MUX2_X1 i_123_0_498 (.A(\o_buffer[87] [13]), .B(i_mem_data[13]), .S(n_32), 
      .Z(n_123_461));
   MUX2_X1 i_123_0_499 (.A(\o_buffer[87] [12]), .B(i_mem_data[12]), .S(n_32), 
      .Z(n_123_460));
   MUX2_X1 i_123_0_500 (.A(\o_buffer[87] [11]), .B(i_mem_data[11]), .S(n_32), 
      .Z(n_123_459));
   MUX2_X1 i_123_0_501 (.A(\o_buffer[87] [10]), .B(i_mem_data[10]), .S(n_32), 
      .Z(n_123_458));
   MUX2_X1 i_123_0_502 (.A(\o_buffer[87] [9]), .B(i_mem_data[9]), .S(n_32), 
      .Z(n_123_457));
   MUX2_X1 i_123_0_503 (.A(\o_buffer[87] [8]), .B(i_mem_data[8]), .S(n_32), 
      .Z(n_123_456));
   MUX2_X1 i_123_0_504 (.A(\o_buffer[87] [7]), .B(i_mem_data[7]), .S(n_32), 
      .Z(n_123_455));
   MUX2_X1 i_123_0_505 (.A(\o_buffer[87] [6]), .B(i_mem_data[6]), .S(n_32), 
      .Z(n_123_454));
   MUX2_X1 i_123_0_506 (.A(\o_buffer[87] [5]), .B(i_mem_data[5]), .S(n_32), 
      .Z(n_123_453));
   MUX2_X1 i_123_0_507 (.A(\o_buffer[87] [4]), .B(i_mem_data[4]), .S(n_32), 
      .Z(n_123_452));
   MUX2_X1 i_123_0_508 (.A(\o_buffer[87] [3]), .B(i_mem_data[3]), .S(n_32), 
      .Z(n_123_451));
   MUX2_X1 i_123_0_509 (.A(\o_buffer[87] [2]), .B(i_mem_data[2]), .S(n_32), 
      .Z(n_123_450));
   MUX2_X1 i_123_0_510 (.A(\o_buffer[87] [1]), .B(i_mem_data[1]), .S(n_32), 
      .Z(n_123_449));
   MUX2_X1 i_123_0_511 (.A(\o_buffer[87] [0]), .B(i_mem_data[0]), .S(n_32), 
      .Z(n_123_448));
   MUX2_X1 i_123_0_512 (.A(\o_buffer[86] [15]), .B(i_mem_data[15]), .S(n_33), 
      .Z(n_123_447));
   MUX2_X1 i_123_0_513 (.A(\o_buffer[86] [14]), .B(i_mem_data[14]), .S(n_33), 
      .Z(n_123_446));
   MUX2_X1 i_123_0_514 (.A(\o_buffer[86] [13]), .B(i_mem_data[13]), .S(n_33), 
      .Z(n_123_445));
   MUX2_X1 i_123_0_515 (.A(\o_buffer[86] [12]), .B(i_mem_data[12]), .S(n_33), 
      .Z(n_123_444));
   MUX2_X1 i_123_0_516 (.A(\o_buffer[86] [11]), .B(i_mem_data[11]), .S(n_33), 
      .Z(n_123_443));
   MUX2_X1 i_123_0_517 (.A(\o_buffer[86] [10]), .B(i_mem_data[10]), .S(n_33), 
      .Z(n_123_442));
   MUX2_X1 i_123_0_518 (.A(\o_buffer[86] [9]), .B(i_mem_data[9]), .S(n_33), 
      .Z(n_123_441));
   MUX2_X1 i_123_0_519 (.A(\o_buffer[86] [8]), .B(i_mem_data[8]), .S(n_33), 
      .Z(n_123_440));
   MUX2_X1 i_123_0_520 (.A(\o_buffer[86] [7]), .B(i_mem_data[7]), .S(n_33), 
      .Z(n_123_439));
   MUX2_X1 i_123_0_521 (.A(\o_buffer[86] [6]), .B(i_mem_data[6]), .S(n_33), 
      .Z(n_123_438));
   MUX2_X1 i_123_0_522 (.A(\o_buffer[86] [5]), .B(i_mem_data[5]), .S(n_33), 
      .Z(n_123_437));
   MUX2_X1 i_123_0_523 (.A(\o_buffer[86] [4]), .B(i_mem_data[4]), .S(n_33), 
      .Z(n_123_436));
   MUX2_X1 i_123_0_524 (.A(\o_buffer[86] [3]), .B(i_mem_data[3]), .S(n_33), 
      .Z(n_123_435));
   MUX2_X1 i_123_0_525 (.A(\o_buffer[86] [2]), .B(i_mem_data[2]), .S(n_33), 
      .Z(n_123_434));
   MUX2_X1 i_123_0_526 (.A(\o_buffer[86] [1]), .B(i_mem_data[1]), .S(n_33), 
      .Z(n_123_433));
   MUX2_X1 i_123_0_527 (.A(\o_buffer[86] [0]), .B(i_mem_data[0]), .S(n_33), 
      .Z(n_123_432));
   MUX2_X1 i_123_0_528 (.A(\o_buffer[85] [15]), .B(i_mem_data[15]), .S(n_34), 
      .Z(n_123_431));
   MUX2_X1 i_123_0_529 (.A(\o_buffer[85] [14]), .B(i_mem_data[14]), .S(n_34), 
      .Z(n_123_430));
   MUX2_X1 i_123_0_530 (.A(\o_buffer[85] [13]), .B(i_mem_data[13]), .S(n_34), 
      .Z(n_123_429));
   MUX2_X1 i_123_0_531 (.A(\o_buffer[85] [12]), .B(i_mem_data[12]), .S(n_34), 
      .Z(n_123_428));
   MUX2_X1 i_123_0_532 (.A(\o_buffer[85] [11]), .B(i_mem_data[11]), .S(n_34), 
      .Z(n_123_427));
   MUX2_X1 i_123_0_533 (.A(\o_buffer[85] [10]), .B(i_mem_data[10]), .S(n_34), 
      .Z(n_123_426));
   MUX2_X1 i_123_0_534 (.A(\o_buffer[85] [9]), .B(i_mem_data[9]), .S(n_34), 
      .Z(n_123_425));
   MUX2_X1 i_123_0_535 (.A(\o_buffer[85] [8]), .B(i_mem_data[8]), .S(n_34), 
      .Z(n_123_424));
   MUX2_X1 i_123_0_536 (.A(\o_buffer[85] [7]), .B(i_mem_data[7]), .S(n_34), 
      .Z(n_123_423));
   MUX2_X1 i_123_0_537 (.A(\o_buffer[85] [6]), .B(i_mem_data[6]), .S(n_34), 
      .Z(n_123_422));
   MUX2_X1 i_123_0_538 (.A(\o_buffer[85] [5]), .B(i_mem_data[5]), .S(n_34), 
      .Z(n_123_421));
   MUX2_X1 i_123_0_539 (.A(\o_buffer[85] [4]), .B(i_mem_data[4]), .S(n_34), 
      .Z(n_123_420));
   MUX2_X1 i_123_0_540 (.A(\o_buffer[85] [3]), .B(i_mem_data[3]), .S(n_34), 
      .Z(n_123_419));
   MUX2_X1 i_123_0_541 (.A(\o_buffer[85] [2]), .B(i_mem_data[2]), .S(n_34), 
      .Z(n_123_418));
   MUX2_X1 i_123_0_542 (.A(\o_buffer[85] [1]), .B(i_mem_data[1]), .S(n_34), 
      .Z(n_123_417));
   MUX2_X1 i_123_0_543 (.A(\o_buffer[85] [0]), .B(i_mem_data[0]), .S(n_34), 
      .Z(n_123_416));
   MUX2_X1 i_123_0_544 (.A(\o_buffer[84] [15]), .B(i_mem_data[15]), .S(n_35), 
      .Z(n_123_415));
   MUX2_X1 i_123_0_545 (.A(\o_buffer[84] [14]), .B(i_mem_data[14]), .S(n_35), 
      .Z(n_123_414));
   MUX2_X1 i_123_0_546 (.A(\o_buffer[84] [13]), .B(i_mem_data[13]), .S(n_35), 
      .Z(n_123_413));
   MUX2_X1 i_123_0_547 (.A(\o_buffer[84] [12]), .B(i_mem_data[12]), .S(n_35), 
      .Z(n_123_412));
   MUX2_X1 i_123_0_548 (.A(\o_buffer[84] [11]), .B(i_mem_data[11]), .S(n_35), 
      .Z(n_123_411));
   MUX2_X1 i_123_0_549 (.A(\o_buffer[84] [10]), .B(i_mem_data[10]), .S(n_35), 
      .Z(n_123_410));
   MUX2_X1 i_123_0_550 (.A(\o_buffer[84] [9]), .B(i_mem_data[9]), .S(n_35), 
      .Z(n_123_409));
   MUX2_X1 i_123_0_551 (.A(\o_buffer[84] [8]), .B(i_mem_data[8]), .S(n_35), 
      .Z(n_123_408));
   MUX2_X1 i_123_0_552 (.A(\o_buffer[84] [7]), .B(i_mem_data[7]), .S(n_35), 
      .Z(n_123_407));
   MUX2_X1 i_123_0_553 (.A(\o_buffer[84] [6]), .B(i_mem_data[6]), .S(n_35), 
      .Z(n_123_406));
   MUX2_X1 i_123_0_554 (.A(\o_buffer[84] [5]), .B(i_mem_data[5]), .S(n_35), 
      .Z(n_123_405));
   MUX2_X1 i_123_0_555 (.A(\o_buffer[84] [4]), .B(i_mem_data[4]), .S(n_35), 
      .Z(n_123_404));
   MUX2_X1 i_123_0_556 (.A(\o_buffer[84] [3]), .B(i_mem_data[3]), .S(n_35), 
      .Z(n_123_403));
   MUX2_X1 i_123_0_557 (.A(\o_buffer[84] [2]), .B(i_mem_data[2]), .S(n_35), 
      .Z(n_123_402));
   MUX2_X1 i_123_0_558 (.A(\o_buffer[84] [1]), .B(i_mem_data[1]), .S(n_35), 
      .Z(n_123_401));
   MUX2_X1 i_123_0_559 (.A(\o_buffer[84] [0]), .B(i_mem_data[0]), .S(n_35), 
      .Z(n_123_400));
   MUX2_X1 i_123_0_560 (.A(\o_buffer[83] [15]), .B(i_mem_data[15]), .S(n_36), 
      .Z(n_123_399));
   MUX2_X1 i_123_0_561 (.A(\o_buffer[83] [14]), .B(i_mem_data[14]), .S(n_36), 
      .Z(n_123_398));
   MUX2_X1 i_123_0_562 (.A(\o_buffer[83] [13]), .B(i_mem_data[13]), .S(n_36), 
      .Z(n_123_397));
   MUX2_X1 i_123_0_563 (.A(\o_buffer[83] [12]), .B(i_mem_data[12]), .S(n_36), 
      .Z(n_123_396));
   MUX2_X1 i_123_0_564 (.A(\o_buffer[83] [11]), .B(i_mem_data[11]), .S(n_36), 
      .Z(n_123_395));
   MUX2_X1 i_123_0_565 (.A(\o_buffer[83] [10]), .B(i_mem_data[10]), .S(n_36), 
      .Z(n_123_394));
   MUX2_X1 i_123_0_566 (.A(\o_buffer[83] [9]), .B(i_mem_data[9]), .S(n_36), 
      .Z(n_123_393));
   MUX2_X1 i_123_0_567 (.A(\o_buffer[83] [8]), .B(i_mem_data[8]), .S(n_36), 
      .Z(n_123_392));
   MUX2_X1 i_123_0_568 (.A(\o_buffer[83] [7]), .B(i_mem_data[7]), .S(n_36), 
      .Z(n_123_391));
   MUX2_X1 i_123_0_569 (.A(\o_buffer[83] [6]), .B(i_mem_data[6]), .S(n_36), 
      .Z(n_123_390));
   MUX2_X1 i_123_0_570 (.A(\o_buffer[83] [5]), .B(i_mem_data[5]), .S(n_36), 
      .Z(n_123_389));
   MUX2_X1 i_123_0_571 (.A(\o_buffer[83] [4]), .B(i_mem_data[4]), .S(n_36), 
      .Z(n_123_388));
   MUX2_X1 i_123_0_572 (.A(\o_buffer[83] [3]), .B(i_mem_data[3]), .S(n_36), 
      .Z(n_123_387));
   MUX2_X1 i_123_0_573 (.A(\o_buffer[83] [2]), .B(i_mem_data[2]), .S(n_36), 
      .Z(n_123_386));
   MUX2_X1 i_123_0_574 (.A(\o_buffer[83] [1]), .B(i_mem_data[1]), .S(n_36), 
      .Z(n_123_385));
   MUX2_X1 i_123_0_575 (.A(\o_buffer[83] [0]), .B(i_mem_data[0]), .S(n_36), 
      .Z(n_123_384));
   MUX2_X1 i_123_0_576 (.A(\o_buffer[82] [15]), .B(i_mem_data[15]), .S(n_37), 
      .Z(n_123_383));
   MUX2_X1 i_123_0_577 (.A(\o_buffer[82] [14]), .B(i_mem_data[14]), .S(n_37), 
      .Z(n_123_382));
   MUX2_X1 i_123_0_578 (.A(\o_buffer[82] [13]), .B(i_mem_data[13]), .S(n_37), 
      .Z(n_123_381));
   MUX2_X1 i_123_0_579 (.A(\o_buffer[82] [12]), .B(i_mem_data[12]), .S(n_37), 
      .Z(n_123_380));
   MUX2_X1 i_123_0_580 (.A(\o_buffer[82] [11]), .B(i_mem_data[11]), .S(n_37), 
      .Z(n_123_379));
   MUX2_X1 i_123_0_581 (.A(\o_buffer[82] [10]), .B(i_mem_data[10]), .S(n_37), 
      .Z(n_123_378));
   MUX2_X1 i_123_0_582 (.A(\o_buffer[82] [9]), .B(i_mem_data[9]), .S(n_37), 
      .Z(n_123_377));
   MUX2_X1 i_123_0_583 (.A(\o_buffer[82] [8]), .B(i_mem_data[8]), .S(n_37), 
      .Z(n_123_376));
   MUX2_X1 i_123_0_584 (.A(\o_buffer[82] [7]), .B(i_mem_data[7]), .S(n_37), 
      .Z(n_123_375));
   MUX2_X1 i_123_0_585 (.A(\o_buffer[82] [6]), .B(i_mem_data[6]), .S(n_37), 
      .Z(n_123_374));
   MUX2_X1 i_123_0_586 (.A(\o_buffer[82] [5]), .B(i_mem_data[5]), .S(n_37), 
      .Z(n_123_373));
   MUX2_X1 i_123_0_587 (.A(\o_buffer[82] [4]), .B(i_mem_data[4]), .S(n_37), 
      .Z(n_123_372));
   MUX2_X1 i_123_0_588 (.A(\o_buffer[82] [3]), .B(i_mem_data[3]), .S(n_37), 
      .Z(n_123_371));
   MUX2_X1 i_123_0_589 (.A(\o_buffer[82] [2]), .B(i_mem_data[2]), .S(n_37), 
      .Z(n_123_370));
   MUX2_X1 i_123_0_590 (.A(\o_buffer[82] [1]), .B(i_mem_data[1]), .S(n_37), 
      .Z(n_123_369));
   MUX2_X1 i_123_0_591 (.A(\o_buffer[82] [0]), .B(i_mem_data[0]), .S(n_37), 
      .Z(n_123_368));
   MUX2_X1 i_123_0_592 (.A(\o_buffer[81] [15]), .B(i_mem_data[15]), .S(n_38), 
      .Z(n_123_367));
   MUX2_X1 i_123_0_593 (.A(\o_buffer[81] [14]), .B(i_mem_data[14]), .S(n_38), 
      .Z(n_123_366));
   MUX2_X1 i_123_0_594 (.A(\o_buffer[81] [13]), .B(i_mem_data[13]), .S(n_38), 
      .Z(n_123_365));
   MUX2_X1 i_123_0_595 (.A(\o_buffer[81] [12]), .B(i_mem_data[12]), .S(n_38), 
      .Z(n_123_364));
   MUX2_X1 i_123_0_596 (.A(\o_buffer[81] [11]), .B(i_mem_data[11]), .S(n_38), 
      .Z(n_123_363));
   MUX2_X1 i_123_0_597 (.A(\o_buffer[81] [10]), .B(i_mem_data[10]), .S(n_38), 
      .Z(n_123_362));
   MUX2_X1 i_123_0_598 (.A(\o_buffer[81] [9]), .B(i_mem_data[9]), .S(n_38), 
      .Z(n_123_361));
   MUX2_X1 i_123_0_599 (.A(\o_buffer[81] [8]), .B(i_mem_data[8]), .S(n_38), 
      .Z(n_123_360));
   MUX2_X1 i_123_0_600 (.A(\o_buffer[81] [7]), .B(i_mem_data[7]), .S(n_38), 
      .Z(n_123_359));
   MUX2_X1 i_123_0_601 (.A(\o_buffer[81] [6]), .B(i_mem_data[6]), .S(n_38), 
      .Z(n_123_358));
   MUX2_X1 i_123_0_602 (.A(\o_buffer[81] [5]), .B(i_mem_data[5]), .S(n_38), 
      .Z(n_123_357));
   MUX2_X1 i_123_0_603 (.A(\o_buffer[81] [4]), .B(i_mem_data[4]), .S(n_38), 
      .Z(n_123_356));
   MUX2_X1 i_123_0_604 (.A(\o_buffer[81] [3]), .B(i_mem_data[3]), .S(n_38), 
      .Z(n_123_355));
   MUX2_X1 i_123_0_605 (.A(\o_buffer[81] [2]), .B(i_mem_data[2]), .S(n_38), 
      .Z(n_123_354));
   MUX2_X1 i_123_0_606 (.A(\o_buffer[81] [1]), .B(i_mem_data[1]), .S(n_38), 
      .Z(n_123_353));
   MUX2_X1 i_123_0_607 (.A(\o_buffer[81] [0]), .B(i_mem_data[0]), .S(n_38), 
      .Z(n_123_352));
   MUX2_X1 i_123_0_608 (.A(\o_buffer[80] [15]), .B(i_mem_data[15]), .S(n_39), 
      .Z(n_123_351));
   MUX2_X1 i_123_0_609 (.A(\o_buffer[80] [14]), .B(i_mem_data[14]), .S(n_39), 
      .Z(n_123_350));
   MUX2_X1 i_123_0_610 (.A(\o_buffer[80] [13]), .B(i_mem_data[13]), .S(n_39), 
      .Z(n_123_349));
   MUX2_X1 i_123_0_611 (.A(\o_buffer[80] [12]), .B(i_mem_data[12]), .S(n_39), 
      .Z(n_123_348));
   MUX2_X1 i_123_0_612 (.A(\o_buffer[80] [11]), .B(i_mem_data[11]), .S(n_39), 
      .Z(n_123_347));
   MUX2_X1 i_123_0_613 (.A(\o_buffer[80] [10]), .B(i_mem_data[10]), .S(n_39), 
      .Z(n_123_346));
   MUX2_X1 i_123_0_614 (.A(\o_buffer[80] [9]), .B(i_mem_data[9]), .S(n_39), 
      .Z(n_123_345));
   MUX2_X1 i_123_0_615 (.A(\o_buffer[80] [8]), .B(i_mem_data[8]), .S(n_39), 
      .Z(n_123_344));
   MUX2_X1 i_123_0_616 (.A(\o_buffer[80] [7]), .B(i_mem_data[7]), .S(n_39), 
      .Z(n_123_343));
   MUX2_X1 i_123_0_617 (.A(\o_buffer[80] [6]), .B(i_mem_data[6]), .S(n_39), 
      .Z(n_123_342));
   MUX2_X1 i_123_0_618 (.A(\o_buffer[80] [5]), .B(i_mem_data[5]), .S(n_39), 
      .Z(n_123_341));
   MUX2_X1 i_123_0_619 (.A(\o_buffer[80] [4]), .B(i_mem_data[4]), .S(n_39), 
      .Z(n_123_340));
   MUX2_X1 i_123_0_620 (.A(\o_buffer[80] [3]), .B(i_mem_data[3]), .S(n_39), 
      .Z(n_123_339));
   MUX2_X1 i_123_0_621 (.A(\o_buffer[80] [2]), .B(i_mem_data[2]), .S(n_39), 
      .Z(n_123_338));
   MUX2_X1 i_123_0_622 (.A(\o_buffer[80] [1]), .B(i_mem_data[1]), .S(n_39), 
      .Z(n_123_337));
   MUX2_X1 i_123_0_623 (.A(\o_buffer[80] [0]), .B(i_mem_data[0]), .S(n_39), 
      .Z(n_123_336));
   MUX2_X1 i_123_0_624 (.A(\o_buffer[79] [15]), .B(i_mem_data[15]), .S(n_40), 
      .Z(n_123_335));
   MUX2_X1 i_123_0_625 (.A(\o_buffer[79] [14]), .B(i_mem_data[14]), .S(n_40), 
      .Z(n_123_334));
   MUX2_X1 i_123_0_626 (.A(\o_buffer[79] [13]), .B(i_mem_data[13]), .S(n_40), 
      .Z(n_123_333));
   MUX2_X1 i_123_0_627 (.A(\o_buffer[79] [12]), .B(i_mem_data[12]), .S(n_40), 
      .Z(n_123_332));
   MUX2_X1 i_123_0_628 (.A(\o_buffer[79] [11]), .B(i_mem_data[11]), .S(n_40), 
      .Z(n_123_331));
   MUX2_X1 i_123_0_629 (.A(\o_buffer[79] [10]), .B(i_mem_data[10]), .S(n_40), 
      .Z(n_123_330));
   MUX2_X1 i_123_0_630 (.A(\o_buffer[79] [9]), .B(i_mem_data[9]), .S(n_40), 
      .Z(n_123_329));
   MUX2_X1 i_123_0_631 (.A(\o_buffer[79] [8]), .B(i_mem_data[8]), .S(n_40), 
      .Z(n_123_328));
   MUX2_X1 i_123_0_632 (.A(\o_buffer[79] [7]), .B(i_mem_data[7]), .S(n_40), 
      .Z(n_123_327));
   MUX2_X1 i_123_0_633 (.A(\o_buffer[79] [6]), .B(i_mem_data[6]), .S(n_40), 
      .Z(n_123_326));
   MUX2_X1 i_123_0_634 (.A(\o_buffer[79] [5]), .B(i_mem_data[5]), .S(n_40), 
      .Z(n_123_325));
   MUX2_X1 i_123_0_635 (.A(\o_buffer[79] [4]), .B(i_mem_data[4]), .S(n_40), 
      .Z(n_123_324));
   MUX2_X1 i_123_0_636 (.A(\o_buffer[79] [3]), .B(i_mem_data[3]), .S(n_40), 
      .Z(n_123_323));
   MUX2_X1 i_123_0_637 (.A(\o_buffer[79] [2]), .B(i_mem_data[2]), .S(n_40), 
      .Z(n_123_322));
   MUX2_X1 i_123_0_638 (.A(\o_buffer[79] [1]), .B(i_mem_data[1]), .S(n_40), 
      .Z(n_123_321));
   MUX2_X1 i_123_0_639 (.A(\o_buffer[79] [0]), .B(i_mem_data[0]), .S(n_40), 
      .Z(n_123_320));
   MUX2_X1 i_123_0_640 (.A(\o_buffer[78] [15]), .B(i_mem_data[15]), .S(n_41), 
      .Z(n_123_319));
   MUX2_X1 i_123_0_641 (.A(\o_buffer[78] [14]), .B(i_mem_data[14]), .S(n_41), 
      .Z(n_123_318));
   MUX2_X1 i_123_0_642 (.A(\o_buffer[78] [13]), .B(i_mem_data[13]), .S(n_41), 
      .Z(n_123_317));
   MUX2_X1 i_123_0_643 (.A(\o_buffer[78] [12]), .B(i_mem_data[12]), .S(n_41), 
      .Z(n_123_316));
   MUX2_X1 i_123_0_644 (.A(\o_buffer[78] [11]), .B(i_mem_data[11]), .S(n_41), 
      .Z(n_123_315));
   MUX2_X1 i_123_0_645 (.A(\o_buffer[78] [10]), .B(i_mem_data[10]), .S(n_41), 
      .Z(n_123_314));
   MUX2_X1 i_123_0_646 (.A(\o_buffer[78] [9]), .B(i_mem_data[9]), .S(n_41), 
      .Z(n_123_313));
   MUX2_X1 i_123_0_647 (.A(\o_buffer[78] [8]), .B(i_mem_data[8]), .S(n_41), 
      .Z(n_123_312));
   MUX2_X1 i_123_0_648 (.A(\o_buffer[78] [7]), .B(i_mem_data[7]), .S(n_41), 
      .Z(n_123_311));
   MUX2_X1 i_123_0_649 (.A(\o_buffer[78] [6]), .B(i_mem_data[6]), .S(n_41), 
      .Z(n_123_310));
   MUX2_X1 i_123_0_650 (.A(\o_buffer[78] [5]), .B(i_mem_data[5]), .S(n_41), 
      .Z(n_123_309));
   MUX2_X1 i_123_0_651 (.A(\o_buffer[78] [4]), .B(i_mem_data[4]), .S(n_41), 
      .Z(n_123_308));
   MUX2_X1 i_123_0_652 (.A(\o_buffer[78] [3]), .B(i_mem_data[3]), .S(n_41), 
      .Z(n_123_307));
   MUX2_X1 i_123_0_653 (.A(\o_buffer[78] [2]), .B(i_mem_data[2]), .S(n_41), 
      .Z(n_123_306));
   MUX2_X1 i_123_0_654 (.A(\o_buffer[78] [1]), .B(i_mem_data[1]), .S(n_41), 
      .Z(n_123_305));
   MUX2_X1 i_123_0_655 (.A(\o_buffer[78] [0]), .B(i_mem_data[0]), .S(n_41), 
      .Z(n_123_304));
   MUX2_X1 i_123_0_656 (.A(\o_buffer[77] [15]), .B(i_mem_data[15]), .S(n_42), 
      .Z(n_123_303));
   MUX2_X1 i_123_0_657 (.A(\o_buffer[77] [14]), .B(i_mem_data[14]), .S(n_42), 
      .Z(n_123_302));
   MUX2_X1 i_123_0_658 (.A(\o_buffer[77] [13]), .B(i_mem_data[13]), .S(n_42), 
      .Z(n_123_301));
   MUX2_X1 i_123_0_659 (.A(\o_buffer[77] [12]), .B(i_mem_data[12]), .S(n_42), 
      .Z(n_123_300));
   MUX2_X1 i_123_0_660 (.A(\o_buffer[77] [11]), .B(i_mem_data[11]), .S(n_42), 
      .Z(n_123_299));
   MUX2_X1 i_123_0_661 (.A(\o_buffer[77] [10]), .B(i_mem_data[10]), .S(n_42), 
      .Z(n_123_298));
   MUX2_X1 i_123_0_662 (.A(\o_buffer[77] [9]), .B(i_mem_data[9]), .S(n_42), 
      .Z(n_123_297));
   MUX2_X1 i_123_0_663 (.A(\o_buffer[77] [8]), .B(i_mem_data[8]), .S(n_42), 
      .Z(n_123_296));
   MUX2_X1 i_123_0_664 (.A(\o_buffer[77] [7]), .B(i_mem_data[7]), .S(n_42), 
      .Z(n_123_295));
   MUX2_X1 i_123_0_665 (.A(\o_buffer[77] [6]), .B(i_mem_data[6]), .S(n_42), 
      .Z(n_123_294));
   MUX2_X1 i_123_0_666 (.A(\o_buffer[77] [5]), .B(i_mem_data[5]), .S(n_42), 
      .Z(n_123_293));
   MUX2_X1 i_123_0_667 (.A(\o_buffer[77] [4]), .B(i_mem_data[4]), .S(n_42), 
      .Z(n_123_292));
   MUX2_X1 i_123_0_668 (.A(\o_buffer[77] [3]), .B(i_mem_data[3]), .S(n_42), 
      .Z(n_123_291));
   MUX2_X1 i_123_0_669 (.A(\o_buffer[77] [2]), .B(i_mem_data[2]), .S(n_42), 
      .Z(n_123_290));
   MUX2_X1 i_123_0_670 (.A(\o_buffer[77] [1]), .B(i_mem_data[1]), .S(n_42), 
      .Z(n_123_289));
   MUX2_X1 i_123_0_671 (.A(\o_buffer[77] [0]), .B(i_mem_data[0]), .S(n_42), 
      .Z(n_123_288));
   MUX2_X1 i_123_0_672 (.A(\o_buffer[76] [15]), .B(i_mem_data[15]), .S(n_43), 
      .Z(n_123_287));
   MUX2_X1 i_123_0_673 (.A(\o_buffer[76] [14]), .B(i_mem_data[14]), .S(n_43), 
      .Z(n_123_286));
   MUX2_X1 i_123_0_674 (.A(\o_buffer[76] [13]), .B(i_mem_data[13]), .S(n_43), 
      .Z(n_123_285));
   MUX2_X1 i_123_0_675 (.A(\o_buffer[76] [12]), .B(i_mem_data[12]), .S(n_43), 
      .Z(n_123_284));
   MUX2_X1 i_123_0_676 (.A(\o_buffer[76] [11]), .B(i_mem_data[11]), .S(n_43), 
      .Z(n_123_283));
   MUX2_X1 i_123_0_677 (.A(\o_buffer[76] [10]), .B(i_mem_data[10]), .S(n_43), 
      .Z(n_123_282));
   MUX2_X1 i_123_0_678 (.A(\o_buffer[76] [9]), .B(i_mem_data[9]), .S(n_43), 
      .Z(n_123_281));
   MUX2_X1 i_123_0_679 (.A(\o_buffer[76] [8]), .B(i_mem_data[8]), .S(n_43), 
      .Z(n_123_280));
   MUX2_X1 i_123_0_680 (.A(\o_buffer[76] [7]), .B(i_mem_data[7]), .S(n_43), 
      .Z(n_123_279));
   MUX2_X1 i_123_0_681 (.A(\o_buffer[76] [6]), .B(i_mem_data[6]), .S(n_43), 
      .Z(n_123_278));
   MUX2_X1 i_123_0_682 (.A(\o_buffer[76] [5]), .B(i_mem_data[5]), .S(n_43), 
      .Z(n_123_277));
   MUX2_X1 i_123_0_683 (.A(\o_buffer[76] [4]), .B(i_mem_data[4]), .S(n_43), 
      .Z(n_123_276));
   MUX2_X1 i_123_0_684 (.A(\o_buffer[76] [3]), .B(i_mem_data[3]), .S(n_43), 
      .Z(n_123_275));
   MUX2_X1 i_123_0_685 (.A(\o_buffer[76] [2]), .B(i_mem_data[2]), .S(n_43), 
      .Z(n_123_274));
   MUX2_X1 i_123_0_686 (.A(\o_buffer[76] [1]), .B(i_mem_data[1]), .S(n_43), 
      .Z(n_123_273));
   MUX2_X1 i_123_0_687 (.A(\o_buffer[76] [0]), .B(i_mem_data[0]), .S(n_43), 
      .Z(n_123_272));
   MUX2_X1 i_123_0_688 (.A(\o_buffer[75] [15]), .B(i_mem_data[15]), .S(n_44), 
      .Z(n_123_271));
   MUX2_X1 i_123_0_689 (.A(\o_buffer[75] [14]), .B(i_mem_data[14]), .S(n_44), 
      .Z(n_123_270));
   MUX2_X1 i_123_0_690 (.A(\o_buffer[75] [13]), .B(i_mem_data[13]), .S(n_44), 
      .Z(n_123_269));
   MUX2_X1 i_123_0_691 (.A(\o_buffer[75] [12]), .B(i_mem_data[12]), .S(n_44), 
      .Z(n_123_268));
   MUX2_X1 i_123_0_692 (.A(\o_buffer[75] [11]), .B(i_mem_data[11]), .S(n_44), 
      .Z(n_123_267));
   MUX2_X1 i_123_0_693 (.A(\o_buffer[75] [10]), .B(i_mem_data[10]), .S(n_44), 
      .Z(n_123_266));
   MUX2_X1 i_123_0_694 (.A(\o_buffer[75] [9]), .B(i_mem_data[9]), .S(n_44), 
      .Z(n_123_265));
   MUX2_X1 i_123_0_695 (.A(\o_buffer[75] [8]), .B(i_mem_data[8]), .S(n_44), 
      .Z(n_123_264));
   MUX2_X1 i_123_0_696 (.A(\o_buffer[75] [7]), .B(i_mem_data[7]), .S(n_44), 
      .Z(n_123_263));
   MUX2_X1 i_123_0_697 (.A(\o_buffer[75] [6]), .B(i_mem_data[6]), .S(n_44), 
      .Z(n_123_262));
   MUX2_X1 i_123_0_698 (.A(\o_buffer[75] [5]), .B(i_mem_data[5]), .S(n_44), 
      .Z(n_123_261));
   MUX2_X1 i_123_0_699 (.A(\o_buffer[75] [4]), .B(i_mem_data[4]), .S(n_44), 
      .Z(n_123_260));
   MUX2_X1 i_123_0_700 (.A(\o_buffer[75] [3]), .B(i_mem_data[3]), .S(n_44), 
      .Z(n_123_259));
   MUX2_X1 i_123_0_701 (.A(\o_buffer[75] [2]), .B(i_mem_data[2]), .S(n_44), 
      .Z(n_123_258));
   MUX2_X1 i_123_0_702 (.A(\o_buffer[75] [1]), .B(i_mem_data[1]), .S(n_44), 
      .Z(n_123_257));
   MUX2_X1 i_123_0_703 (.A(\o_buffer[75] [0]), .B(i_mem_data[0]), .S(n_44), 
      .Z(n_123_256));
   MUX2_X1 i_123_0_704 (.A(\o_buffer[74] [15]), .B(i_mem_data[15]), .S(n_45), 
      .Z(n_123_255));
   MUX2_X1 i_123_0_705 (.A(\o_buffer[74] [14]), .B(i_mem_data[14]), .S(n_45), 
      .Z(n_123_254));
   MUX2_X1 i_123_0_706 (.A(\o_buffer[74] [13]), .B(i_mem_data[13]), .S(n_45), 
      .Z(n_123_253));
   MUX2_X1 i_123_0_707 (.A(\o_buffer[74] [12]), .B(i_mem_data[12]), .S(n_45), 
      .Z(n_123_252));
   MUX2_X1 i_123_0_708 (.A(\o_buffer[74] [11]), .B(i_mem_data[11]), .S(n_45), 
      .Z(n_123_251));
   MUX2_X1 i_123_0_709 (.A(\o_buffer[74] [10]), .B(i_mem_data[10]), .S(n_45), 
      .Z(n_123_250));
   MUX2_X1 i_123_0_710 (.A(\o_buffer[74] [9]), .B(i_mem_data[9]), .S(n_45), 
      .Z(n_123_249));
   MUX2_X1 i_123_0_711 (.A(\o_buffer[74] [8]), .B(i_mem_data[8]), .S(n_45), 
      .Z(n_123_248));
   MUX2_X1 i_123_0_712 (.A(\o_buffer[74] [7]), .B(i_mem_data[7]), .S(n_45), 
      .Z(n_123_247));
   MUX2_X1 i_123_0_713 (.A(\o_buffer[74] [6]), .B(i_mem_data[6]), .S(n_45), 
      .Z(n_123_246));
   MUX2_X1 i_123_0_714 (.A(\o_buffer[74] [5]), .B(i_mem_data[5]), .S(n_45), 
      .Z(n_123_245));
   MUX2_X1 i_123_0_715 (.A(\o_buffer[74] [4]), .B(i_mem_data[4]), .S(n_45), 
      .Z(n_123_244));
   MUX2_X1 i_123_0_716 (.A(\o_buffer[74] [3]), .B(i_mem_data[3]), .S(n_45), 
      .Z(n_123_243));
   MUX2_X1 i_123_0_717 (.A(\o_buffer[74] [2]), .B(i_mem_data[2]), .S(n_45), 
      .Z(n_123_242));
   MUX2_X1 i_123_0_718 (.A(\o_buffer[74] [1]), .B(i_mem_data[1]), .S(n_45), 
      .Z(n_123_241));
   MUX2_X1 i_123_0_719 (.A(\o_buffer[74] [0]), .B(i_mem_data[0]), .S(n_45), 
      .Z(n_123_240));
   MUX2_X1 i_123_0_720 (.A(\o_buffer[73] [15]), .B(i_mem_data[15]), .S(n_46), 
      .Z(n_123_239));
   MUX2_X1 i_123_0_721 (.A(\o_buffer[73] [14]), .B(i_mem_data[14]), .S(n_46), 
      .Z(n_123_238));
   MUX2_X1 i_123_0_722 (.A(\o_buffer[73] [13]), .B(i_mem_data[13]), .S(n_46), 
      .Z(n_123_237));
   MUX2_X1 i_123_0_723 (.A(\o_buffer[73] [12]), .B(i_mem_data[12]), .S(n_46), 
      .Z(n_123_236));
   MUX2_X1 i_123_0_724 (.A(\o_buffer[73] [11]), .B(i_mem_data[11]), .S(n_46), 
      .Z(n_123_235));
   MUX2_X1 i_123_0_725 (.A(\o_buffer[73] [10]), .B(i_mem_data[10]), .S(n_46), 
      .Z(n_123_234));
   MUX2_X1 i_123_0_726 (.A(\o_buffer[73] [9]), .B(i_mem_data[9]), .S(n_46), 
      .Z(n_123_233));
   MUX2_X1 i_123_0_727 (.A(\o_buffer[73] [8]), .B(i_mem_data[8]), .S(n_46), 
      .Z(n_123_232));
   MUX2_X1 i_123_0_728 (.A(\o_buffer[73] [7]), .B(i_mem_data[7]), .S(n_46), 
      .Z(n_123_231));
   MUX2_X1 i_123_0_729 (.A(\o_buffer[73] [6]), .B(i_mem_data[6]), .S(n_46), 
      .Z(n_123_230));
   MUX2_X1 i_123_0_730 (.A(\o_buffer[73] [5]), .B(i_mem_data[5]), .S(n_46), 
      .Z(n_123_229));
   MUX2_X1 i_123_0_731 (.A(\o_buffer[73] [4]), .B(i_mem_data[4]), .S(n_46), 
      .Z(n_123_228));
   MUX2_X1 i_123_0_732 (.A(\o_buffer[73] [3]), .B(i_mem_data[3]), .S(n_46), 
      .Z(n_123_227));
   MUX2_X1 i_123_0_733 (.A(\o_buffer[73] [2]), .B(i_mem_data[2]), .S(n_46), 
      .Z(n_123_226));
   MUX2_X1 i_123_0_734 (.A(\o_buffer[73] [1]), .B(i_mem_data[1]), .S(n_46), 
      .Z(n_123_225));
   MUX2_X1 i_123_0_735 (.A(\o_buffer[73] [0]), .B(i_mem_data[0]), .S(n_46), 
      .Z(n_123_224));
   MUX2_X1 i_123_0_736 (.A(\o_buffer[72] [15]), .B(i_mem_data[15]), .S(n_47), 
      .Z(n_123_223));
   MUX2_X1 i_123_0_737 (.A(\o_buffer[72] [14]), .B(i_mem_data[14]), .S(n_47), 
      .Z(n_123_222));
   MUX2_X1 i_123_0_738 (.A(\o_buffer[72] [13]), .B(i_mem_data[13]), .S(n_47), 
      .Z(n_123_221));
   MUX2_X1 i_123_0_739 (.A(\o_buffer[72] [12]), .B(i_mem_data[12]), .S(n_47), 
      .Z(n_123_220));
   MUX2_X1 i_123_0_740 (.A(\o_buffer[72] [11]), .B(i_mem_data[11]), .S(n_47), 
      .Z(n_123_219));
   MUX2_X1 i_123_0_741 (.A(\o_buffer[72] [10]), .B(i_mem_data[10]), .S(n_47), 
      .Z(n_123_218));
   MUX2_X1 i_123_0_742 (.A(\o_buffer[72] [9]), .B(i_mem_data[9]), .S(n_47), 
      .Z(n_123_217));
   MUX2_X1 i_123_0_743 (.A(\o_buffer[72] [8]), .B(i_mem_data[8]), .S(n_47), 
      .Z(n_123_216));
   MUX2_X1 i_123_0_744 (.A(\o_buffer[72] [7]), .B(i_mem_data[7]), .S(n_47), 
      .Z(n_123_215));
   MUX2_X1 i_123_0_745 (.A(\o_buffer[72] [6]), .B(i_mem_data[6]), .S(n_47), 
      .Z(n_123_214));
   MUX2_X1 i_123_0_746 (.A(\o_buffer[72] [5]), .B(i_mem_data[5]), .S(n_47), 
      .Z(n_123_213));
   MUX2_X1 i_123_0_747 (.A(\o_buffer[72] [4]), .B(i_mem_data[4]), .S(n_47), 
      .Z(n_123_212));
   MUX2_X1 i_123_0_748 (.A(\o_buffer[72] [3]), .B(i_mem_data[3]), .S(n_47), 
      .Z(n_123_211));
   MUX2_X1 i_123_0_749 (.A(\o_buffer[72] [2]), .B(i_mem_data[2]), .S(n_47), 
      .Z(n_123_210));
   MUX2_X1 i_123_0_750 (.A(\o_buffer[72] [1]), .B(i_mem_data[1]), .S(n_47), 
      .Z(n_123_209));
   MUX2_X1 i_123_0_751 (.A(\o_buffer[72] [0]), .B(i_mem_data[0]), .S(n_47), 
      .Z(n_123_208));
   MUX2_X1 i_123_0_752 (.A(\o_buffer[71] [15]), .B(i_mem_data[15]), .S(n_48), 
      .Z(n_123_207));
   MUX2_X1 i_123_0_753 (.A(\o_buffer[71] [14]), .B(i_mem_data[14]), .S(n_48), 
      .Z(n_123_206));
   MUX2_X1 i_123_0_754 (.A(\o_buffer[71] [13]), .B(i_mem_data[13]), .S(n_48), 
      .Z(n_123_205));
   MUX2_X1 i_123_0_755 (.A(\o_buffer[71] [12]), .B(i_mem_data[12]), .S(n_48), 
      .Z(n_123_204));
   MUX2_X1 i_123_0_756 (.A(\o_buffer[71] [11]), .B(i_mem_data[11]), .S(n_48), 
      .Z(n_123_203));
   MUX2_X1 i_123_0_757 (.A(\o_buffer[71] [10]), .B(i_mem_data[10]), .S(n_48), 
      .Z(n_123_202));
   MUX2_X1 i_123_0_758 (.A(\o_buffer[71] [9]), .B(i_mem_data[9]), .S(n_48), 
      .Z(n_123_201));
   MUX2_X1 i_123_0_759 (.A(\o_buffer[71] [8]), .B(i_mem_data[8]), .S(n_48), 
      .Z(n_123_200));
   MUX2_X1 i_123_0_760 (.A(\o_buffer[71] [7]), .B(i_mem_data[7]), .S(n_48), 
      .Z(n_123_199));
   MUX2_X1 i_123_0_761 (.A(\o_buffer[71] [6]), .B(i_mem_data[6]), .S(n_48), 
      .Z(n_123_198));
   MUX2_X1 i_123_0_762 (.A(\o_buffer[71] [5]), .B(i_mem_data[5]), .S(n_48), 
      .Z(n_123_197));
   MUX2_X1 i_123_0_763 (.A(\o_buffer[71] [4]), .B(i_mem_data[4]), .S(n_48), 
      .Z(n_123_196));
   MUX2_X1 i_123_0_764 (.A(\o_buffer[71] [3]), .B(i_mem_data[3]), .S(n_48), 
      .Z(n_123_195));
   MUX2_X1 i_123_0_765 (.A(\o_buffer[71] [2]), .B(i_mem_data[2]), .S(n_48), 
      .Z(n_123_194));
   MUX2_X1 i_123_0_766 (.A(\o_buffer[71] [1]), .B(i_mem_data[1]), .S(n_48), 
      .Z(n_123_193));
   MUX2_X1 i_123_0_767 (.A(\o_buffer[71] [0]), .B(i_mem_data[0]), .S(n_48), 
      .Z(n_123_192));
   MUX2_X1 i_123_0_768 (.A(\o_buffer[70] [15]), .B(i_mem_data[15]), .S(n_49), 
      .Z(n_123_191));
   MUX2_X1 i_123_0_769 (.A(\o_buffer[70] [14]), .B(i_mem_data[14]), .S(n_49), 
      .Z(n_123_190));
   MUX2_X1 i_123_0_770 (.A(\o_buffer[70] [13]), .B(i_mem_data[13]), .S(n_49), 
      .Z(n_123_189));
   MUX2_X1 i_123_0_771 (.A(\o_buffer[70] [12]), .B(i_mem_data[12]), .S(n_49), 
      .Z(n_123_188));
   MUX2_X1 i_123_0_772 (.A(\o_buffer[70] [11]), .B(i_mem_data[11]), .S(n_49), 
      .Z(n_123_187));
   MUX2_X1 i_123_0_773 (.A(\o_buffer[70] [10]), .B(i_mem_data[10]), .S(n_49), 
      .Z(n_123_186));
   MUX2_X1 i_123_0_774 (.A(\o_buffer[70] [9]), .B(i_mem_data[9]), .S(n_49), 
      .Z(n_123_185));
   MUX2_X1 i_123_0_775 (.A(\o_buffer[70] [8]), .B(i_mem_data[8]), .S(n_49), 
      .Z(n_123_184));
   MUX2_X1 i_123_0_776 (.A(\o_buffer[70] [7]), .B(i_mem_data[7]), .S(n_49), 
      .Z(n_123_183));
   MUX2_X1 i_123_0_777 (.A(\o_buffer[70] [6]), .B(i_mem_data[6]), .S(n_49), 
      .Z(n_123_182));
   MUX2_X1 i_123_0_778 (.A(\o_buffer[70] [5]), .B(i_mem_data[5]), .S(n_49), 
      .Z(n_123_181));
   MUX2_X1 i_123_0_779 (.A(\o_buffer[70] [4]), .B(i_mem_data[4]), .S(n_49), 
      .Z(n_123_180));
   MUX2_X1 i_123_0_780 (.A(\o_buffer[70] [3]), .B(i_mem_data[3]), .S(n_49), 
      .Z(n_123_179));
   MUX2_X1 i_123_0_781 (.A(\o_buffer[70] [2]), .B(i_mem_data[2]), .S(n_49), 
      .Z(n_123_178));
   MUX2_X1 i_123_0_782 (.A(\o_buffer[70] [1]), .B(i_mem_data[1]), .S(n_49), 
      .Z(n_123_177));
   MUX2_X1 i_123_0_783 (.A(\o_buffer[70] [0]), .B(i_mem_data[0]), .S(n_49), 
      .Z(n_123_176));
   MUX2_X1 i_123_0_784 (.A(\o_buffer[69] [15]), .B(i_mem_data[15]), .S(n_50), 
      .Z(n_123_175));
   MUX2_X1 i_123_0_785 (.A(\o_buffer[69] [14]), .B(i_mem_data[14]), .S(n_50), 
      .Z(n_123_174));
   MUX2_X1 i_123_0_786 (.A(\o_buffer[69] [13]), .B(i_mem_data[13]), .S(n_50), 
      .Z(n_123_173));
   MUX2_X1 i_123_0_787 (.A(\o_buffer[69] [12]), .B(i_mem_data[12]), .S(n_50), 
      .Z(n_123_172));
   MUX2_X1 i_123_0_788 (.A(\o_buffer[69] [11]), .B(i_mem_data[11]), .S(n_50), 
      .Z(n_123_171));
   MUX2_X1 i_123_0_789 (.A(\o_buffer[69] [10]), .B(i_mem_data[10]), .S(n_50), 
      .Z(n_123_170));
   MUX2_X1 i_123_0_790 (.A(\o_buffer[69] [9]), .B(i_mem_data[9]), .S(n_50), 
      .Z(n_123_169));
   MUX2_X1 i_123_0_791 (.A(\o_buffer[69] [8]), .B(i_mem_data[8]), .S(n_50), 
      .Z(n_123_168));
   MUX2_X1 i_123_0_792 (.A(\o_buffer[69] [7]), .B(i_mem_data[7]), .S(n_50), 
      .Z(n_123_167));
   MUX2_X1 i_123_0_793 (.A(\o_buffer[69] [6]), .B(i_mem_data[6]), .S(n_50), 
      .Z(n_123_166));
   MUX2_X1 i_123_0_794 (.A(\o_buffer[69] [5]), .B(i_mem_data[5]), .S(n_50), 
      .Z(n_123_165));
   MUX2_X1 i_123_0_795 (.A(\o_buffer[69] [4]), .B(i_mem_data[4]), .S(n_50), 
      .Z(n_123_164));
   MUX2_X1 i_123_0_796 (.A(\o_buffer[69] [3]), .B(i_mem_data[3]), .S(n_50), 
      .Z(n_123_163));
   MUX2_X1 i_123_0_797 (.A(\o_buffer[69] [2]), .B(i_mem_data[2]), .S(n_50), 
      .Z(n_123_162));
   MUX2_X1 i_123_0_798 (.A(\o_buffer[69] [1]), .B(i_mem_data[1]), .S(n_50), 
      .Z(n_123_161));
   MUX2_X1 i_123_0_799 (.A(\o_buffer[69] [0]), .B(i_mem_data[0]), .S(n_50), 
      .Z(n_123_160));
   MUX2_X1 i_123_0_800 (.A(\o_buffer[68] [15]), .B(i_mem_data[15]), .S(n_51), 
      .Z(n_123_159));
   MUX2_X1 i_123_0_801 (.A(\o_buffer[68] [14]), .B(i_mem_data[14]), .S(n_51), 
      .Z(n_123_158));
   MUX2_X1 i_123_0_802 (.A(\o_buffer[68] [13]), .B(i_mem_data[13]), .S(n_51), 
      .Z(n_123_157));
   MUX2_X1 i_123_0_803 (.A(\o_buffer[68] [12]), .B(i_mem_data[12]), .S(n_51), 
      .Z(n_123_156));
   MUX2_X1 i_123_0_804 (.A(\o_buffer[68] [11]), .B(i_mem_data[11]), .S(n_51), 
      .Z(n_123_155));
   MUX2_X1 i_123_0_805 (.A(\o_buffer[68] [10]), .B(i_mem_data[10]), .S(n_51), 
      .Z(n_123_154));
   MUX2_X1 i_123_0_806 (.A(\o_buffer[68] [9]), .B(i_mem_data[9]), .S(n_51), 
      .Z(n_123_153));
   MUX2_X1 i_123_0_807 (.A(\o_buffer[68] [8]), .B(i_mem_data[8]), .S(n_51), 
      .Z(n_123_152));
   MUX2_X1 i_123_0_808 (.A(\o_buffer[68] [7]), .B(i_mem_data[7]), .S(n_51), 
      .Z(n_123_151));
   MUX2_X1 i_123_0_809 (.A(\o_buffer[68] [6]), .B(i_mem_data[6]), .S(n_51), 
      .Z(n_123_150));
   MUX2_X1 i_123_0_810 (.A(\o_buffer[68] [5]), .B(i_mem_data[5]), .S(n_51), 
      .Z(n_123_149));
   MUX2_X1 i_123_0_811 (.A(\o_buffer[68] [4]), .B(i_mem_data[4]), .S(n_51), 
      .Z(n_123_148));
   MUX2_X1 i_123_0_812 (.A(\o_buffer[68] [3]), .B(i_mem_data[3]), .S(n_51), 
      .Z(n_123_147));
   MUX2_X1 i_123_0_813 (.A(\o_buffer[68] [2]), .B(i_mem_data[2]), .S(n_51), 
      .Z(n_123_146));
   MUX2_X1 i_123_0_814 (.A(\o_buffer[68] [1]), .B(i_mem_data[1]), .S(n_51), 
      .Z(n_123_145));
   MUX2_X1 i_123_0_815 (.A(\o_buffer[68] [0]), .B(i_mem_data[0]), .S(n_51), 
      .Z(n_123_144));
   MUX2_X1 i_123_0_816 (.A(\o_buffer[67] [15]), .B(i_mem_data[15]), .S(n_52), 
      .Z(n_123_143));
   MUX2_X1 i_123_0_817 (.A(\o_buffer[67] [14]), .B(i_mem_data[14]), .S(n_52), 
      .Z(n_123_142));
   MUX2_X1 i_123_0_818 (.A(\o_buffer[67] [13]), .B(i_mem_data[13]), .S(n_52), 
      .Z(n_123_141));
   MUX2_X1 i_123_0_819 (.A(\o_buffer[67] [12]), .B(i_mem_data[12]), .S(n_52), 
      .Z(n_123_140));
   MUX2_X1 i_123_0_820 (.A(\o_buffer[67] [11]), .B(i_mem_data[11]), .S(n_52), 
      .Z(n_123_139));
   MUX2_X1 i_123_0_821 (.A(\o_buffer[67] [10]), .B(i_mem_data[10]), .S(n_52), 
      .Z(n_123_138));
   MUX2_X1 i_123_0_822 (.A(\o_buffer[67] [9]), .B(i_mem_data[9]), .S(n_52), 
      .Z(n_123_137));
   MUX2_X1 i_123_0_823 (.A(\o_buffer[67] [8]), .B(i_mem_data[8]), .S(n_52), 
      .Z(n_123_136));
   MUX2_X1 i_123_0_824 (.A(\o_buffer[67] [7]), .B(i_mem_data[7]), .S(n_52), 
      .Z(n_123_135));
   MUX2_X1 i_123_0_825 (.A(\o_buffer[67] [6]), .B(i_mem_data[6]), .S(n_52), 
      .Z(n_123_134));
   MUX2_X1 i_123_0_826 (.A(\o_buffer[67] [5]), .B(i_mem_data[5]), .S(n_52), 
      .Z(n_123_133));
   MUX2_X1 i_123_0_827 (.A(\o_buffer[67] [4]), .B(i_mem_data[4]), .S(n_52), 
      .Z(n_123_132));
   MUX2_X1 i_123_0_828 (.A(\o_buffer[67] [3]), .B(i_mem_data[3]), .S(n_52), 
      .Z(n_123_131));
   MUX2_X1 i_123_0_829 (.A(\o_buffer[67] [2]), .B(i_mem_data[2]), .S(n_52), 
      .Z(n_123_130));
   MUX2_X1 i_123_0_830 (.A(\o_buffer[67] [1]), .B(i_mem_data[1]), .S(n_52), 
      .Z(n_123_129));
   MUX2_X1 i_123_0_831 (.A(\o_buffer[67] [0]), .B(i_mem_data[0]), .S(n_52), 
      .Z(n_123_128));
   MUX2_X1 i_123_0_832 (.A(\o_buffer[66] [15]), .B(i_mem_data[15]), .S(n_53), 
      .Z(n_123_127));
   MUX2_X1 i_123_0_833 (.A(\o_buffer[66] [14]), .B(i_mem_data[14]), .S(n_53), 
      .Z(n_123_126));
   MUX2_X1 i_123_0_834 (.A(\o_buffer[66] [13]), .B(i_mem_data[13]), .S(n_53), 
      .Z(n_123_125));
   MUX2_X1 i_123_0_835 (.A(\o_buffer[66] [12]), .B(i_mem_data[12]), .S(n_53), 
      .Z(n_123_124));
   MUX2_X1 i_123_0_836 (.A(\o_buffer[66] [11]), .B(i_mem_data[11]), .S(n_53), 
      .Z(n_123_123));
   MUX2_X1 i_123_0_837 (.A(\o_buffer[66] [10]), .B(i_mem_data[10]), .S(n_53), 
      .Z(n_123_122));
   MUX2_X1 i_123_0_838 (.A(\o_buffer[66] [9]), .B(i_mem_data[9]), .S(n_53), 
      .Z(n_123_121));
   MUX2_X1 i_123_0_839 (.A(\o_buffer[66] [8]), .B(i_mem_data[8]), .S(n_53), 
      .Z(n_123_120));
   MUX2_X1 i_123_0_840 (.A(\o_buffer[66] [7]), .B(i_mem_data[7]), .S(n_53), 
      .Z(n_123_119));
   MUX2_X1 i_123_0_841 (.A(\o_buffer[66] [6]), .B(i_mem_data[6]), .S(n_53), 
      .Z(n_123_118));
   MUX2_X1 i_123_0_842 (.A(\o_buffer[66] [5]), .B(i_mem_data[5]), .S(n_53), 
      .Z(n_123_117));
   MUX2_X1 i_123_0_843 (.A(\o_buffer[66] [4]), .B(i_mem_data[4]), .S(n_53), 
      .Z(n_123_116));
   MUX2_X1 i_123_0_844 (.A(\o_buffer[66] [3]), .B(i_mem_data[3]), .S(n_53), 
      .Z(n_123_115));
   MUX2_X1 i_123_0_845 (.A(\o_buffer[66] [2]), .B(i_mem_data[2]), .S(n_53), 
      .Z(n_123_114));
   MUX2_X1 i_123_0_846 (.A(\o_buffer[66] [1]), .B(i_mem_data[1]), .S(n_53), 
      .Z(n_123_113));
   MUX2_X1 i_123_0_847 (.A(\o_buffer[66] [0]), .B(i_mem_data[0]), .S(n_53), 
      .Z(n_123_112));
   MUX2_X1 i_123_0_848 (.A(\o_buffer[65] [15]), .B(i_mem_data[15]), .S(n_54), 
      .Z(n_123_111));
   MUX2_X1 i_123_0_849 (.A(\o_buffer[65] [14]), .B(i_mem_data[14]), .S(n_54), 
      .Z(n_123_110));
   MUX2_X1 i_123_0_850 (.A(\o_buffer[65] [13]), .B(i_mem_data[13]), .S(n_54), 
      .Z(n_123_109));
   MUX2_X1 i_123_0_851 (.A(\o_buffer[65] [12]), .B(i_mem_data[12]), .S(n_54), 
      .Z(n_123_108));
   MUX2_X1 i_123_0_852 (.A(\o_buffer[65] [11]), .B(i_mem_data[11]), .S(n_54), 
      .Z(n_123_107));
   MUX2_X1 i_123_0_853 (.A(\o_buffer[65] [10]), .B(i_mem_data[10]), .S(n_54), 
      .Z(n_123_106));
   MUX2_X1 i_123_0_854 (.A(\o_buffer[65] [9]), .B(i_mem_data[9]), .S(n_54), 
      .Z(n_123_105));
   MUX2_X1 i_123_0_855 (.A(\o_buffer[65] [8]), .B(i_mem_data[8]), .S(n_54), 
      .Z(n_123_104));
   MUX2_X1 i_123_0_856 (.A(\o_buffer[65] [7]), .B(i_mem_data[7]), .S(n_54), 
      .Z(n_123_103));
   MUX2_X1 i_123_0_857 (.A(\o_buffer[65] [6]), .B(i_mem_data[6]), .S(n_54), 
      .Z(n_123_102));
   MUX2_X1 i_123_0_858 (.A(\o_buffer[65] [5]), .B(i_mem_data[5]), .S(n_54), 
      .Z(n_123_101));
   MUX2_X1 i_123_0_859 (.A(\o_buffer[65] [4]), .B(i_mem_data[4]), .S(n_54), 
      .Z(n_123_100));
   MUX2_X1 i_123_0_860 (.A(\o_buffer[65] [3]), .B(i_mem_data[3]), .S(n_54), 
      .Z(n_123_99));
   MUX2_X1 i_123_0_861 (.A(\o_buffer[65] [2]), .B(i_mem_data[2]), .S(n_54), 
      .Z(n_123_98));
   MUX2_X1 i_123_0_862 (.A(\o_buffer[65] [1]), .B(i_mem_data[1]), .S(n_54), 
      .Z(n_123_97));
   MUX2_X1 i_123_0_863 (.A(\o_buffer[65] [0]), .B(i_mem_data[0]), .S(n_54), 
      .Z(n_123_96));
   MUX2_X1 i_123_0_864 (.A(\o_buffer[64] [15]), .B(i_mem_data[15]), .S(n_55), 
      .Z(n_123_95));
   MUX2_X1 i_123_0_865 (.A(\o_buffer[64] [14]), .B(i_mem_data[14]), .S(n_55), 
      .Z(n_123_94));
   MUX2_X1 i_123_0_866 (.A(\o_buffer[64] [13]), .B(i_mem_data[13]), .S(n_55), 
      .Z(n_123_93));
   MUX2_X1 i_123_0_867 (.A(\o_buffer[64] [12]), .B(i_mem_data[12]), .S(n_55), 
      .Z(n_123_92));
   MUX2_X1 i_123_0_868 (.A(\o_buffer[64] [11]), .B(i_mem_data[11]), .S(n_55), 
      .Z(n_123_91));
   MUX2_X1 i_123_0_869 (.A(\o_buffer[64] [10]), .B(i_mem_data[10]), .S(n_55), 
      .Z(n_123_90));
   MUX2_X1 i_123_0_870 (.A(\o_buffer[64] [9]), .B(i_mem_data[9]), .S(n_55), 
      .Z(n_123_89));
   MUX2_X1 i_123_0_871 (.A(\o_buffer[64] [8]), .B(i_mem_data[8]), .S(n_55), 
      .Z(n_123_88));
   MUX2_X1 i_123_0_872 (.A(\o_buffer[64] [7]), .B(i_mem_data[7]), .S(n_55), 
      .Z(n_123_87));
   MUX2_X1 i_123_0_873 (.A(\o_buffer[64] [6]), .B(i_mem_data[6]), .S(n_55), 
      .Z(n_123_86));
   MUX2_X1 i_123_0_874 (.A(\o_buffer[64] [5]), .B(i_mem_data[5]), .S(n_55), 
      .Z(n_123_85));
   MUX2_X1 i_123_0_875 (.A(\o_buffer[64] [4]), .B(i_mem_data[4]), .S(n_55), 
      .Z(n_123_84));
   MUX2_X1 i_123_0_876 (.A(\o_buffer[64] [3]), .B(i_mem_data[3]), .S(n_55), 
      .Z(n_123_83));
   MUX2_X1 i_123_0_877 (.A(\o_buffer[64] [2]), .B(i_mem_data[2]), .S(n_55), 
      .Z(n_123_82));
   MUX2_X1 i_123_0_878 (.A(\o_buffer[64] [1]), .B(i_mem_data[1]), .S(n_55), 
      .Z(n_123_81));
   MUX2_X1 i_123_0_879 (.A(\o_buffer[64] [0]), .B(i_mem_data[0]), .S(n_55), 
      .Z(n_123_80));
   MUX2_X1 i_123_0_880 (.A(\o_buffer[63] [15]), .B(i_mem_data[15]), .S(n_56), 
      .Z(n_123_79));
   MUX2_X1 i_123_0_881 (.A(\o_buffer[63] [14]), .B(i_mem_data[14]), .S(n_56), 
      .Z(n_123_78));
   MUX2_X1 i_123_0_882 (.A(\o_buffer[63] [13]), .B(i_mem_data[13]), .S(n_56), 
      .Z(n_123_77));
   MUX2_X1 i_123_0_883 (.A(\o_buffer[63] [12]), .B(i_mem_data[12]), .S(n_56), 
      .Z(n_123_76));
   MUX2_X1 i_123_0_884 (.A(\o_buffer[63] [11]), .B(i_mem_data[11]), .S(n_56), 
      .Z(n_123_75));
   MUX2_X1 i_123_0_885 (.A(\o_buffer[63] [10]), .B(i_mem_data[10]), .S(n_56), 
      .Z(n_123_74));
   MUX2_X1 i_123_0_886 (.A(\o_buffer[63] [9]), .B(i_mem_data[9]), .S(n_56), 
      .Z(n_123_73));
   MUX2_X1 i_123_0_887 (.A(\o_buffer[63] [8]), .B(i_mem_data[8]), .S(n_56), 
      .Z(n_123_72));
   MUX2_X1 i_123_0_888 (.A(\o_buffer[63] [7]), .B(i_mem_data[7]), .S(n_56), 
      .Z(n_123_71));
   MUX2_X1 i_123_0_889 (.A(\o_buffer[63] [6]), .B(i_mem_data[6]), .S(n_56), 
      .Z(n_123_70));
   MUX2_X1 i_123_0_890 (.A(\o_buffer[63] [5]), .B(i_mem_data[5]), .S(n_56), 
      .Z(n_123_69));
   MUX2_X1 i_123_0_891 (.A(\o_buffer[63] [4]), .B(i_mem_data[4]), .S(n_56), 
      .Z(n_123_68));
   MUX2_X1 i_123_0_892 (.A(\o_buffer[63] [3]), .B(i_mem_data[3]), .S(n_56), 
      .Z(n_123_67));
   MUX2_X1 i_123_0_893 (.A(\o_buffer[63] [2]), .B(i_mem_data[2]), .S(n_56), 
      .Z(n_123_66));
   MUX2_X1 i_123_0_894 (.A(\o_buffer[63] [1]), .B(i_mem_data[1]), .S(n_56), 
      .Z(n_123_65));
   MUX2_X1 i_123_0_895 (.A(\o_buffer[63] [0]), .B(i_mem_data[0]), .S(n_56), 
      .Z(n_123_64));
   MUX2_X1 i_123_0_896 (.A(\o_buffer[62] [15]), .B(i_mem_data[15]), .S(n_57), 
      .Z(n_123_63));
   MUX2_X1 i_123_0_897 (.A(\o_buffer[62] [14]), .B(i_mem_data[14]), .S(n_57), 
      .Z(n_123_62));
   MUX2_X1 i_123_0_898 (.A(\o_buffer[62] [13]), .B(i_mem_data[13]), .S(n_57), 
      .Z(n_123_61));
   MUX2_X1 i_123_0_899 (.A(\o_buffer[62] [12]), .B(i_mem_data[12]), .S(n_57), 
      .Z(n_123_60));
   MUX2_X1 i_123_0_900 (.A(\o_buffer[62] [11]), .B(i_mem_data[11]), .S(n_57), 
      .Z(n_123_59));
   MUX2_X1 i_123_0_901 (.A(\o_buffer[62] [10]), .B(i_mem_data[10]), .S(n_57), 
      .Z(n_123_58));
   MUX2_X1 i_123_0_902 (.A(\o_buffer[62] [9]), .B(i_mem_data[9]), .S(n_57), 
      .Z(n_123_57));
   MUX2_X1 i_123_0_903 (.A(\o_buffer[62] [8]), .B(i_mem_data[8]), .S(n_57), 
      .Z(n_123_56));
   MUX2_X1 i_123_0_904 (.A(\o_buffer[62] [7]), .B(i_mem_data[7]), .S(n_57), 
      .Z(n_123_55));
   MUX2_X1 i_123_0_905 (.A(\o_buffer[62] [6]), .B(i_mem_data[6]), .S(n_57), 
      .Z(n_123_54));
   MUX2_X1 i_123_0_906 (.A(\o_buffer[62] [5]), .B(i_mem_data[5]), .S(n_57), 
      .Z(n_123_53));
   MUX2_X1 i_123_0_907 (.A(\o_buffer[62] [4]), .B(i_mem_data[4]), .S(n_57), 
      .Z(n_123_52));
   MUX2_X1 i_123_0_908 (.A(\o_buffer[62] [3]), .B(i_mem_data[3]), .S(n_57), 
      .Z(n_123_51));
   MUX2_X1 i_123_0_909 (.A(\o_buffer[62] [2]), .B(i_mem_data[2]), .S(n_57), 
      .Z(n_123_50));
   MUX2_X1 i_123_0_910 (.A(\o_buffer[62] [1]), .B(i_mem_data[1]), .S(n_57), 
      .Z(n_123_49));
   MUX2_X1 i_123_0_911 (.A(\o_buffer[62] [0]), .B(i_mem_data[0]), .S(n_57), 
      .Z(n_123_48));
   MUX2_X1 i_123_0_912 (.A(\o_buffer[61] [15]), .B(i_mem_data[15]), .S(n_58), 
      .Z(n_123_47));
   MUX2_X1 i_123_0_913 (.A(\o_buffer[61] [14]), .B(i_mem_data[14]), .S(n_58), 
      .Z(n_123_46));
   MUX2_X1 i_123_0_914 (.A(\o_buffer[61] [13]), .B(i_mem_data[13]), .S(n_58), 
      .Z(n_123_45));
   MUX2_X1 i_123_0_915 (.A(\o_buffer[61] [12]), .B(i_mem_data[12]), .S(n_58), 
      .Z(n_123_44));
   MUX2_X1 i_123_0_916 (.A(\o_buffer[61] [11]), .B(i_mem_data[11]), .S(n_58), 
      .Z(n_123_43));
   MUX2_X1 i_123_0_917 (.A(\o_buffer[61] [10]), .B(i_mem_data[10]), .S(n_58), 
      .Z(n_123_42));
   MUX2_X1 i_123_0_918 (.A(\o_buffer[61] [9]), .B(i_mem_data[9]), .S(n_58), 
      .Z(n_123_41));
   MUX2_X1 i_123_0_919 (.A(\o_buffer[61] [8]), .B(i_mem_data[8]), .S(n_58), 
      .Z(n_123_40));
   MUX2_X1 i_123_0_920 (.A(\o_buffer[61] [7]), .B(i_mem_data[7]), .S(n_58), 
      .Z(n_123_39));
   MUX2_X1 i_123_0_921 (.A(\o_buffer[61] [6]), .B(i_mem_data[6]), .S(n_58), 
      .Z(n_123_38));
   MUX2_X1 i_123_0_922 (.A(\o_buffer[61] [5]), .B(i_mem_data[5]), .S(n_58), 
      .Z(n_123_37));
   MUX2_X1 i_123_0_923 (.A(\o_buffer[61] [4]), .B(i_mem_data[4]), .S(n_58), 
      .Z(n_123_36));
   MUX2_X1 i_123_0_924 (.A(\o_buffer[61] [3]), .B(i_mem_data[3]), .S(n_58), 
      .Z(n_123_35));
   MUX2_X1 i_123_0_925 (.A(\o_buffer[61] [2]), .B(i_mem_data[2]), .S(n_58), 
      .Z(n_123_34));
   MUX2_X1 i_123_0_926 (.A(\o_buffer[61] [1]), .B(i_mem_data[1]), .S(n_58), 
      .Z(n_123_33));
   MUX2_X1 i_123_0_927 (.A(\o_buffer[61] [0]), .B(i_mem_data[0]), .S(n_58), 
      .Z(n_123_32));
   MUX2_X1 i_123_0_928 (.A(\o_buffer[60] [15]), .B(i_mem_data[15]), .S(n_59), 
      .Z(n_123_31));
   MUX2_X1 i_123_0_929 (.A(\o_buffer[60] [14]), .B(i_mem_data[14]), .S(n_59), 
      .Z(n_123_30));
   MUX2_X1 i_123_0_930 (.A(\o_buffer[60] [13]), .B(i_mem_data[13]), .S(n_59), 
      .Z(n_123_29));
   MUX2_X1 i_123_0_931 (.A(\o_buffer[60] [12]), .B(i_mem_data[12]), .S(n_59), 
      .Z(n_123_28));
   MUX2_X1 i_123_0_932 (.A(\o_buffer[60] [11]), .B(i_mem_data[11]), .S(n_59), 
      .Z(n_123_27));
   MUX2_X1 i_123_0_933 (.A(\o_buffer[60] [10]), .B(i_mem_data[10]), .S(n_59), 
      .Z(n_123_26));
   MUX2_X1 i_123_0_934 (.A(\o_buffer[60] [9]), .B(i_mem_data[9]), .S(n_59), 
      .Z(n_123_25));
   MUX2_X1 i_123_0_935 (.A(\o_buffer[60] [8]), .B(i_mem_data[8]), .S(n_59), 
      .Z(n_123_24));
   MUX2_X1 i_123_0_936 (.A(\o_buffer[60] [7]), .B(i_mem_data[7]), .S(n_59), 
      .Z(n_123_23));
   MUX2_X1 i_123_0_937 (.A(\o_buffer[60] [6]), .B(i_mem_data[6]), .S(n_59), 
      .Z(n_123_22));
   MUX2_X1 i_123_0_938 (.A(\o_buffer[60] [5]), .B(i_mem_data[5]), .S(n_59), 
      .Z(n_123_21));
   MUX2_X1 i_123_0_939 (.A(\o_buffer[60] [4]), .B(i_mem_data[4]), .S(n_59), 
      .Z(n_123_20));
   MUX2_X1 i_123_0_940 (.A(\o_buffer[60] [3]), .B(i_mem_data[3]), .S(n_59), 
      .Z(n_123_19));
   MUX2_X1 i_123_0_941 (.A(\o_buffer[60] [2]), .B(i_mem_data[2]), .S(n_59), 
      .Z(n_123_18));
   MUX2_X1 i_123_0_942 (.A(\o_buffer[60] [1]), .B(i_mem_data[1]), .S(n_59), 
      .Z(n_123_17));
   MUX2_X1 i_123_0_943 (.A(\o_buffer[60] [0]), .B(i_mem_data[0]), .S(n_59), 
      .Z(n_123_16));
   MUX2_X1 i_123_0_944 (.A(\o_buffer[59] [15]), .B(i_mem_data[15]), .S(n_60), 
      .Z(n_123_15));
   MUX2_X1 i_123_0_945 (.A(\o_buffer[59] [14]), .B(i_mem_data[14]), .S(n_60), 
      .Z(n_123_14));
   MUX2_X1 i_123_0_946 (.A(\o_buffer[59] [13]), .B(i_mem_data[13]), .S(n_60), 
      .Z(n_123_13));
   MUX2_X1 i_123_0_947 (.A(\o_buffer[59] [12]), .B(i_mem_data[12]), .S(n_60), 
      .Z(n_123_12));
   MUX2_X1 i_123_0_948 (.A(\o_buffer[59] [11]), .B(i_mem_data[11]), .S(n_60), 
      .Z(n_123_11));
   MUX2_X1 i_123_0_949 (.A(\o_buffer[59] [10]), .B(i_mem_data[10]), .S(n_60), 
      .Z(n_123_10));
   MUX2_X1 i_123_0_950 (.A(\o_buffer[59] [9]), .B(i_mem_data[9]), .S(n_60), 
      .Z(n_123_9));
   MUX2_X1 i_123_0_951 (.A(\o_buffer[59] [8]), .B(i_mem_data[8]), .S(n_60), 
      .Z(n_123_8));
   MUX2_X1 i_123_0_952 (.A(\o_buffer[59] [7]), .B(i_mem_data[7]), .S(n_60), 
      .Z(n_123_7));
   MUX2_X1 i_123_0_953 (.A(\o_buffer[59] [6]), .B(i_mem_data[6]), .S(n_60), 
      .Z(n_123_6));
   MUX2_X1 i_123_0_954 (.A(\o_buffer[59] [5]), .B(i_mem_data[5]), .S(n_60), 
      .Z(n_123_5));
   MUX2_X1 i_123_0_955 (.A(\o_buffer[59] [4]), .B(i_mem_data[4]), .S(n_60), 
      .Z(n_123_4));
   MUX2_X1 i_123_0_956 (.A(\o_buffer[59] [3]), .B(i_mem_data[3]), .S(n_60), 
      .Z(n_123_3));
   MUX2_X1 i_123_0_957 (.A(\o_buffer[59] [2]), .B(i_mem_data[2]), .S(n_60), 
      .Z(n_123_2));
   MUX2_X1 i_123_0_958 (.A(\o_buffer[59] [1]), .B(i_mem_data[1]), .S(n_60), 
      .Z(n_123_1));
   MUX2_X1 i_123_0_959 (.A(\o_buffer[59] [0]), .B(i_mem_data[0]), .S(n_60), 
      .Z(n_123_0));
   DFF_X1 \o_buffer_reg[58][15]  (.D(n_132_959), .CK(n_120), .Q(
      \o_buffer[58] [15]), .QN());
   DFF_X1 \o_buffer_reg[58][14]  (.D(n_132_958), .CK(n_120), .Q(
      \o_buffer[58] [14]), .QN());
   DFF_X1 \o_buffer_reg[58][13]  (.D(n_132_957), .CK(n_120), .Q(
      \o_buffer[58] [13]), .QN());
   DFF_X1 \o_buffer_reg[58][12]  (.D(n_132_956), .CK(n_120), .Q(
      \o_buffer[58] [12]), .QN());
   DFF_X1 \o_buffer_reg[58][11]  (.D(n_132_955), .CK(n_120), .Q(
      \o_buffer[58] [11]), .QN());
   DFF_X1 \o_buffer_reg[58][10]  (.D(n_132_954), .CK(n_120), .Q(
      \o_buffer[58] [10]), .QN());
   DFF_X1 \o_buffer_reg[58][9]  (.D(n_132_953), .CK(n_120), .Q(\o_buffer[58] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][8]  (.D(n_132_952), .CK(n_120), .Q(\o_buffer[58] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][7]  (.D(n_132_951), .CK(n_120), .Q(\o_buffer[58] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][6]  (.D(n_132_950), .CK(n_120), .Q(\o_buffer[58] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][5]  (.D(n_132_949), .CK(n_120), .Q(\o_buffer[58] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][4]  (.D(n_132_948), .CK(n_120), .Q(\o_buffer[58] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][3]  (.D(n_132_947), .CK(n_120), .Q(\o_buffer[58] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][2]  (.D(n_132_946), .CK(n_120), .Q(\o_buffer[58] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][1]  (.D(n_132_945), .CK(n_120), .Q(\o_buffer[58] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[58][0]  (.D(n_132_944), .CK(n_120), .Q(\o_buffer[58] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][15]  (.D(n_132_943), .CK(n_120), .Q(
      \o_buffer[57] [15]), .QN());
   DFF_X1 \o_buffer_reg[57][14]  (.D(n_132_942), .CK(n_120), .Q(
      \o_buffer[57] [14]), .QN());
   DFF_X1 \o_buffer_reg[57][13]  (.D(n_132_941), .CK(n_120), .Q(
      \o_buffer[57] [13]), .QN());
   DFF_X1 \o_buffer_reg[57][12]  (.D(n_132_940), .CK(n_120), .Q(
      \o_buffer[57] [12]), .QN());
   DFF_X1 \o_buffer_reg[57][11]  (.D(n_132_939), .CK(n_120), .Q(
      \o_buffer[57] [11]), .QN());
   DFF_X1 \o_buffer_reg[57][10]  (.D(n_132_938), .CK(n_120), .Q(
      \o_buffer[57] [10]), .QN());
   DFF_X1 \o_buffer_reg[57][9]  (.D(n_132_937), .CK(n_120), .Q(\o_buffer[57] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][8]  (.D(n_132_936), .CK(n_120), .Q(\o_buffer[57] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][7]  (.D(n_132_935), .CK(n_120), .Q(\o_buffer[57] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][6]  (.D(n_132_934), .CK(n_120), .Q(\o_buffer[57] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][5]  (.D(n_132_933), .CK(n_120), .Q(\o_buffer[57] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][4]  (.D(n_132_932), .CK(n_120), .Q(\o_buffer[57] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][3]  (.D(n_132_931), .CK(n_120), .Q(\o_buffer[57] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][2]  (.D(n_132_930), .CK(n_120), .Q(\o_buffer[57] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][1]  (.D(n_132_929), .CK(n_120), .Q(\o_buffer[57] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[57][0]  (.D(n_132_928), .CK(n_120), .Q(\o_buffer[57] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][15]  (.D(n_132_927), .CK(n_120), .Q(
      \o_buffer[56] [15]), .QN());
   DFF_X1 \o_buffer_reg[56][14]  (.D(n_132_926), .CK(n_120), .Q(
      \o_buffer[56] [14]), .QN());
   DFF_X1 \o_buffer_reg[56][13]  (.D(n_132_925), .CK(n_120), .Q(
      \o_buffer[56] [13]), .QN());
   DFF_X1 \o_buffer_reg[56][12]  (.D(n_132_924), .CK(n_120), .Q(
      \o_buffer[56] [12]), .QN());
   DFF_X1 \o_buffer_reg[56][11]  (.D(n_132_923), .CK(n_120), .Q(
      \o_buffer[56] [11]), .QN());
   DFF_X1 \o_buffer_reg[56][10]  (.D(n_132_922), .CK(n_120), .Q(
      \o_buffer[56] [10]), .QN());
   DFF_X1 \o_buffer_reg[56][9]  (.D(n_132_921), .CK(n_120), .Q(\o_buffer[56] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][8]  (.D(n_132_920), .CK(n_120), .Q(\o_buffer[56] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][7]  (.D(n_132_919), .CK(n_120), .Q(\o_buffer[56] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][6]  (.D(n_132_918), .CK(n_120), .Q(\o_buffer[56] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][5]  (.D(n_132_917), .CK(n_120), .Q(\o_buffer[56] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][4]  (.D(n_132_916), .CK(n_120), .Q(\o_buffer[56] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][3]  (.D(n_132_915), .CK(n_120), .Q(\o_buffer[56] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][2]  (.D(n_132_914), .CK(n_120), .Q(\o_buffer[56] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][1]  (.D(n_132_913), .CK(n_120), .Q(\o_buffer[56] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[56][0]  (.D(n_132_912), .CK(n_120), .Q(\o_buffer[56] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][15]  (.D(n_132_911), .CK(n_120), .Q(
      \o_buffer[55] [15]), .QN());
   DFF_X1 \o_buffer_reg[55][14]  (.D(n_132_910), .CK(n_120), .Q(
      \o_buffer[55] [14]), .QN());
   DFF_X1 \o_buffer_reg[55][13]  (.D(n_132_909), .CK(n_120), .Q(
      \o_buffer[55] [13]), .QN());
   DFF_X1 \o_buffer_reg[55][12]  (.D(n_132_908), .CK(n_120), .Q(
      \o_buffer[55] [12]), .QN());
   DFF_X1 \o_buffer_reg[55][11]  (.D(n_132_907), .CK(n_120), .Q(
      \o_buffer[55] [11]), .QN());
   DFF_X1 \o_buffer_reg[55][10]  (.D(n_132_906), .CK(n_120), .Q(
      \o_buffer[55] [10]), .QN());
   DFF_X1 \o_buffer_reg[55][9]  (.D(n_132_905), .CK(n_120), .Q(\o_buffer[55] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][8]  (.D(n_132_904), .CK(n_120), .Q(\o_buffer[55] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][7]  (.D(n_132_903), .CK(n_120), .Q(\o_buffer[55] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][6]  (.D(n_132_902), .CK(n_120), .Q(\o_buffer[55] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][5]  (.D(n_132_901), .CK(n_120), .Q(\o_buffer[55] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][4]  (.D(n_132_900), .CK(n_120), .Q(\o_buffer[55] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][3]  (.D(n_132_899), .CK(n_120), .Q(\o_buffer[55] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][2]  (.D(n_132_898), .CK(n_120), .Q(\o_buffer[55] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][1]  (.D(n_132_897), .CK(n_120), .Q(\o_buffer[55] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[55][0]  (.D(n_132_896), .CK(n_120), .Q(\o_buffer[55] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][15]  (.D(n_132_895), .CK(n_120), .Q(
      \o_buffer[54] [15]), .QN());
   DFF_X1 \o_buffer_reg[54][14]  (.D(n_132_894), .CK(n_120), .Q(
      \o_buffer[54] [14]), .QN());
   DFF_X1 \o_buffer_reg[54][13]  (.D(n_132_893), .CK(n_120), .Q(
      \o_buffer[54] [13]), .QN());
   DFF_X1 \o_buffer_reg[54][12]  (.D(n_132_892), .CK(n_120), .Q(
      \o_buffer[54] [12]), .QN());
   DFF_X1 \o_buffer_reg[54][11]  (.D(n_132_891), .CK(n_120), .Q(
      \o_buffer[54] [11]), .QN());
   DFF_X1 \o_buffer_reg[54][10]  (.D(n_132_890), .CK(n_120), .Q(
      \o_buffer[54] [10]), .QN());
   DFF_X1 \o_buffer_reg[54][9]  (.D(n_132_889), .CK(n_120), .Q(\o_buffer[54] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][8]  (.D(n_132_888), .CK(n_120), .Q(\o_buffer[54] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][7]  (.D(n_132_887), .CK(n_120), .Q(\o_buffer[54] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][6]  (.D(n_132_886), .CK(n_120), .Q(\o_buffer[54] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][5]  (.D(n_132_885), .CK(n_120), .Q(\o_buffer[54] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][4]  (.D(n_132_884), .CK(n_120), .Q(\o_buffer[54] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][3]  (.D(n_132_883), .CK(n_120), .Q(\o_buffer[54] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][2]  (.D(n_132_882), .CK(n_120), .Q(\o_buffer[54] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][1]  (.D(n_132_881), .CK(n_120), .Q(\o_buffer[54] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[54][0]  (.D(n_132_880), .CK(n_120), .Q(\o_buffer[54] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][15]  (.D(n_132_879), .CK(n_120), .Q(
      \o_buffer[53] [15]), .QN());
   DFF_X1 \o_buffer_reg[53][14]  (.D(n_132_878), .CK(n_120), .Q(
      \o_buffer[53] [14]), .QN());
   DFF_X1 \o_buffer_reg[53][13]  (.D(n_132_877), .CK(n_120), .Q(
      \o_buffer[53] [13]), .QN());
   DFF_X1 \o_buffer_reg[53][12]  (.D(n_132_876), .CK(n_120), .Q(
      \o_buffer[53] [12]), .QN());
   DFF_X1 \o_buffer_reg[53][11]  (.D(n_132_875), .CK(n_120), .Q(
      \o_buffer[53] [11]), .QN());
   DFF_X1 \o_buffer_reg[53][10]  (.D(n_132_874), .CK(n_120), .Q(
      \o_buffer[53] [10]), .QN());
   DFF_X1 \o_buffer_reg[53][9]  (.D(n_132_873), .CK(n_120), .Q(\o_buffer[53] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][8]  (.D(n_132_872), .CK(n_120), .Q(\o_buffer[53] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][7]  (.D(n_132_871), .CK(n_120), .Q(\o_buffer[53] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][6]  (.D(n_132_870), .CK(n_120), .Q(\o_buffer[53] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][5]  (.D(n_132_869), .CK(n_120), .Q(\o_buffer[53] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][4]  (.D(n_132_868), .CK(n_120), .Q(\o_buffer[53] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][3]  (.D(n_132_867), .CK(n_120), .Q(\o_buffer[53] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][2]  (.D(n_132_866), .CK(n_120), .Q(\o_buffer[53] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][1]  (.D(n_132_865), .CK(n_120), .Q(\o_buffer[53] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[53][0]  (.D(n_132_864), .CK(n_120), .Q(\o_buffer[53] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][15]  (.D(n_132_863), .CK(n_120), .Q(
      \o_buffer[52] [15]), .QN());
   DFF_X1 \o_buffer_reg[52][14]  (.D(n_132_862), .CK(n_120), .Q(
      \o_buffer[52] [14]), .QN());
   DFF_X1 \o_buffer_reg[52][13]  (.D(n_132_861), .CK(n_120), .Q(
      \o_buffer[52] [13]), .QN());
   DFF_X1 \o_buffer_reg[52][12]  (.D(n_132_860), .CK(n_120), .Q(
      \o_buffer[52] [12]), .QN());
   DFF_X1 \o_buffer_reg[52][11]  (.D(n_132_859), .CK(n_120), .Q(
      \o_buffer[52] [11]), .QN());
   DFF_X1 \o_buffer_reg[52][10]  (.D(n_132_858), .CK(n_120), .Q(
      \o_buffer[52] [10]), .QN());
   DFF_X1 \o_buffer_reg[52][9]  (.D(n_132_857), .CK(n_120), .Q(\o_buffer[52] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][8]  (.D(n_132_856), .CK(n_120), .Q(\o_buffer[52] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][7]  (.D(n_132_855), .CK(n_120), .Q(\o_buffer[52] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][6]  (.D(n_132_854), .CK(n_120), .Q(\o_buffer[52] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][5]  (.D(n_132_853), .CK(n_120), .Q(\o_buffer[52] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][4]  (.D(n_132_852), .CK(n_120), .Q(\o_buffer[52] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][3]  (.D(n_132_851), .CK(n_120), .Q(\o_buffer[52] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][2]  (.D(n_132_850), .CK(n_120), .Q(\o_buffer[52] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][1]  (.D(n_132_849), .CK(n_120), .Q(\o_buffer[52] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[52][0]  (.D(n_132_848), .CK(n_120), .Q(\o_buffer[52] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][15]  (.D(n_132_847), .CK(n_120), .Q(
      \o_buffer[51] [15]), .QN());
   DFF_X1 \o_buffer_reg[51][14]  (.D(n_132_846), .CK(n_120), .Q(
      \o_buffer[51] [14]), .QN());
   DFF_X1 \o_buffer_reg[51][13]  (.D(n_132_845), .CK(n_120), .Q(
      \o_buffer[51] [13]), .QN());
   DFF_X1 \o_buffer_reg[51][12]  (.D(n_132_844), .CK(n_120), .Q(
      \o_buffer[51] [12]), .QN());
   DFF_X1 \o_buffer_reg[51][11]  (.D(n_132_843), .CK(n_120), .Q(
      \o_buffer[51] [11]), .QN());
   DFF_X1 \o_buffer_reg[51][10]  (.D(n_132_842), .CK(n_120), .Q(
      \o_buffer[51] [10]), .QN());
   DFF_X1 \o_buffer_reg[51][9]  (.D(n_132_841), .CK(n_120), .Q(\o_buffer[51] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][8]  (.D(n_132_840), .CK(n_120), .Q(\o_buffer[51] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][7]  (.D(n_132_839), .CK(n_120), .Q(\o_buffer[51] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][6]  (.D(n_132_838), .CK(n_120), .Q(\o_buffer[51] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][5]  (.D(n_132_837), .CK(n_120), .Q(\o_buffer[51] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][4]  (.D(n_132_836), .CK(n_120), .Q(\o_buffer[51] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][3]  (.D(n_132_835), .CK(n_120), .Q(\o_buffer[51] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][2]  (.D(n_132_834), .CK(n_120), .Q(\o_buffer[51] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][1]  (.D(n_132_833), .CK(n_120), .Q(\o_buffer[51] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[51][0]  (.D(n_132_832), .CK(n_120), .Q(\o_buffer[51] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][15]  (.D(n_132_831), .CK(n_120), .Q(
      \o_buffer[50] [15]), .QN());
   DFF_X1 \o_buffer_reg[50][14]  (.D(n_132_830), .CK(n_120), .Q(
      \o_buffer[50] [14]), .QN());
   DFF_X1 \o_buffer_reg[50][13]  (.D(n_132_829), .CK(n_120), .Q(
      \o_buffer[50] [13]), .QN());
   DFF_X1 \o_buffer_reg[50][12]  (.D(n_132_828), .CK(n_120), .Q(
      \o_buffer[50] [12]), .QN());
   DFF_X1 \o_buffer_reg[50][11]  (.D(n_132_827), .CK(n_120), .Q(
      \o_buffer[50] [11]), .QN());
   DFF_X1 \o_buffer_reg[50][10]  (.D(n_132_826), .CK(n_120), .Q(
      \o_buffer[50] [10]), .QN());
   DFF_X1 \o_buffer_reg[50][9]  (.D(n_132_825), .CK(n_120), .Q(\o_buffer[50] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][8]  (.D(n_132_824), .CK(n_120), .Q(\o_buffer[50] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][7]  (.D(n_132_823), .CK(n_120), .Q(\o_buffer[50] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][6]  (.D(n_132_822), .CK(n_120), .Q(\o_buffer[50] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][5]  (.D(n_132_821), .CK(n_120), .Q(\o_buffer[50] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][4]  (.D(n_132_820), .CK(n_120), .Q(\o_buffer[50] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][3]  (.D(n_132_819), .CK(n_120), .Q(\o_buffer[50] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][2]  (.D(n_132_818), .CK(n_120), .Q(\o_buffer[50] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][1]  (.D(n_132_817), .CK(n_120), .Q(\o_buffer[50] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[50][0]  (.D(n_132_816), .CK(n_120), .Q(\o_buffer[50] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][15]  (.D(n_132_815), .CK(n_120), .Q(
      \o_buffer[49] [15]), .QN());
   DFF_X1 \o_buffer_reg[49][14]  (.D(n_132_814), .CK(n_120), .Q(
      \o_buffer[49] [14]), .QN());
   DFF_X1 \o_buffer_reg[49][13]  (.D(n_132_813), .CK(n_120), .Q(
      \o_buffer[49] [13]), .QN());
   DFF_X1 \o_buffer_reg[49][12]  (.D(n_132_812), .CK(n_120), .Q(
      \o_buffer[49] [12]), .QN());
   DFF_X1 \o_buffer_reg[49][11]  (.D(n_132_811), .CK(n_120), .Q(
      \o_buffer[49] [11]), .QN());
   DFF_X1 \o_buffer_reg[49][10]  (.D(n_132_810), .CK(n_120), .Q(
      \o_buffer[49] [10]), .QN());
   DFF_X1 \o_buffer_reg[49][9]  (.D(n_132_809), .CK(n_120), .Q(\o_buffer[49] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][8]  (.D(n_132_808), .CK(n_120), .Q(\o_buffer[49] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][7]  (.D(n_132_807), .CK(n_120), .Q(\o_buffer[49] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][6]  (.D(n_132_806), .CK(n_120), .Q(\o_buffer[49] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][5]  (.D(n_132_805), .CK(n_120), .Q(\o_buffer[49] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][4]  (.D(n_132_804), .CK(n_120), .Q(\o_buffer[49] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][3]  (.D(n_132_803), .CK(n_120), .Q(\o_buffer[49] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][2]  (.D(n_132_802), .CK(n_120), .Q(\o_buffer[49] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][1]  (.D(n_132_801), .CK(n_120), .Q(\o_buffer[49] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[49][0]  (.D(n_132_800), .CK(n_120), .Q(\o_buffer[49] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][15]  (.D(n_132_799), .CK(n_120), .Q(
      \o_buffer[48] [15]), .QN());
   DFF_X1 \o_buffer_reg[48][14]  (.D(n_132_798), .CK(n_120), .Q(
      \o_buffer[48] [14]), .QN());
   DFF_X1 \o_buffer_reg[48][13]  (.D(n_132_797), .CK(n_120), .Q(
      \o_buffer[48] [13]), .QN());
   DFF_X1 \o_buffer_reg[48][12]  (.D(n_132_796), .CK(n_120), .Q(
      \o_buffer[48] [12]), .QN());
   DFF_X1 \o_buffer_reg[48][11]  (.D(n_132_795), .CK(n_120), .Q(
      \o_buffer[48] [11]), .QN());
   DFF_X1 \o_buffer_reg[48][10]  (.D(n_132_794), .CK(n_120), .Q(
      \o_buffer[48] [10]), .QN());
   DFF_X1 \o_buffer_reg[48][9]  (.D(n_132_793), .CK(n_120), .Q(\o_buffer[48] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][8]  (.D(n_132_792), .CK(n_120), .Q(\o_buffer[48] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][7]  (.D(n_132_791), .CK(n_120), .Q(\o_buffer[48] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][6]  (.D(n_132_790), .CK(n_120), .Q(\o_buffer[48] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][5]  (.D(n_132_789), .CK(n_120), .Q(\o_buffer[48] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][4]  (.D(n_132_788), .CK(n_120), .Q(\o_buffer[48] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][3]  (.D(n_132_787), .CK(n_120), .Q(\o_buffer[48] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][2]  (.D(n_132_786), .CK(n_120), .Q(\o_buffer[48] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][1]  (.D(n_132_785), .CK(n_120), .Q(\o_buffer[48] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[48][0]  (.D(n_132_784), .CK(n_120), .Q(\o_buffer[48] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][15]  (.D(n_132_783), .CK(n_120), .Q(
      \o_buffer[47] [15]), .QN());
   DFF_X1 \o_buffer_reg[47][14]  (.D(n_132_782), .CK(n_120), .Q(
      \o_buffer[47] [14]), .QN());
   DFF_X1 \o_buffer_reg[47][13]  (.D(n_132_781), .CK(n_120), .Q(
      \o_buffer[47] [13]), .QN());
   DFF_X1 \o_buffer_reg[47][12]  (.D(n_132_780), .CK(n_120), .Q(
      \o_buffer[47] [12]), .QN());
   DFF_X1 \o_buffer_reg[47][11]  (.D(n_132_779), .CK(n_120), .Q(
      \o_buffer[47] [11]), .QN());
   DFF_X1 \o_buffer_reg[47][10]  (.D(n_132_778), .CK(n_120), .Q(
      \o_buffer[47] [10]), .QN());
   DFF_X1 \o_buffer_reg[47][9]  (.D(n_132_777), .CK(n_120), .Q(\o_buffer[47] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][8]  (.D(n_132_776), .CK(n_120), .Q(\o_buffer[47] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][7]  (.D(n_132_775), .CK(n_120), .Q(\o_buffer[47] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][6]  (.D(n_132_774), .CK(n_120), .Q(\o_buffer[47] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][5]  (.D(n_132_773), .CK(n_120), .Q(\o_buffer[47] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][4]  (.D(n_132_772), .CK(n_120), .Q(\o_buffer[47] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][3]  (.D(n_132_771), .CK(n_120), .Q(\o_buffer[47] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][2]  (.D(n_132_770), .CK(n_120), .Q(\o_buffer[47] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][1]  (.D(n_132_769), .CK(n_120), .Q(\o_buffer[47] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[47][0]  (.D(n_132_768), .CK(n_120), .Q(\o_buffer[47] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][15]  (.D(n_132_767), .CK(n_120), .Q(
      \o_buffer[46] [15]), .QN());
   DFF_X1 \o_buffer_reg[46][14]  (.D(n_132_766), .CK(n_120), .Q(
      \o_buffer[46] [14]), .QN());
   DFF_X1 \o_buffer_reg[46][13]  (.D(n_132_765), .CK(n_120), .Q(
      \o_buffer[46] [13]), .QN());
   DFF_X1 \o_buffer_reg[46][12]  (.D(n_132_764), .CK(n_120), .Q(
      \o_buffer[46] [12]), .QN());
   DFF_X1 \o_buffer_reg[46][11]  (.D(n_132_763), .CK(n_120), .Q(
      \o_buffer[46] [11]), .QN());
   DFF_X1 \o_buffer_reg[46][10]  (.D(n_132_762), .CK(n_120), .Q(
      \o_buffer[46] [10]), .QN());
   DFF_X1 \o_buffer_reg[46][9]  (.D(n_132_761), .CK(n_120), .Q(\o_buffer[46] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][8]  (.D(n_132_760), .CK(n_120), .Q(\o_buffer[46] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][7]  (.D(n_132_759), .CK(n_120), .Q(\o_buffer[46] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][6]  (.D(n_132_758), .CK(n_120), .Q(\o_buffer[46] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][5]  (.D(n_132_757), .CK(n_120), .Q(\o_buffer[46] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][4]  (.D(n_132_756), .CK(n_120), .Q(\o_buffer[46] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][3]  (.D(n_132_755), .CK(n_120), .Q(\o_buffer[46] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][2]  (.D(n_132_754), .CK(n_120), .Q(\o_buffer[46] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][1]  (.D(n_132_753), .CK(n_120), .Q(\o_buffer[46] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[46][0]  (.D(n_132_752), .CK(n_120), .Q(\o_buffer[46] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][15]  (.D(n_132_751), .CK(n_120), .Q(
      \o_buffer[45] [15]), .QN());
   DFF_X1 \o_buffer_reg[45][14]  (.D(n_132_750), .CK(n_120), .Q(
      \o_buffer[45] [14]), .QN());
   DFF_X1 \o_buffer_reg[45][13]  (.D(n_132_749), .CK(n_120), .Q(
      \o_buffer[45] [13]), .QN());
   DFF_X1 \o_buffer_reg[45][12]  (.D(n_132_748), .CK(n_120), .Q(
      \o_buffer[45] [12]), .QN());
   DFF_X1 \o_buffer_reg[45][11]  (.D(n_132_747), .CK(n_120), .Q(
      \o_buffer[45] [11]), .QN());
   DFF_X1 \o_buffer_reg[45][10]  (.D(n_132_746), .CK(n_120), .Q(
      \o_buffer[45] [10]), .QN());
   DFF_X1 \o_buffer_reg[45][9]  (.D(n_132_745), .CK(n_120), .Q(\o_buffer[45] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][8]  (.D(n_132_744), .CK(n_120), .Q(\o_buffer[45] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][7]  (.D(n_132_743), .CK(n_120), .Q(\o_buffer[45] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][6]  (.D(n_132_742), .CK(n_120), .Q(\o_buffer[45] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][5]  (.D(n_132_741), .CK(n_120), .Q(\o_buffer[45] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][4]  (.D(n_132_740), .CK(n_120), .Q(\o_buffer[45] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][3]  (.D(n_132_739), .CK(n_120), .Q(\o_buffer[45] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][2]  (.D(n_132_738), .CK(n_120), .Q(\o_buffer[45] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][1]  (.D(n_132_737), .CK(n_120), .Q(\o_buffer[45] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[45][0]  (.D(n_132_736), .CK(n_120), .Q(\o_buffer[45] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][15]  (.D(n_132_735), .CK(n_120), .Q(
      \o_buffer[44] [15]), .QN());
   DFF_X1 \o_buffer_reg[44][14]  (.D(n_132_734), .CK(n_120), .Q(
      \o_buffer[44] [14]), .QN());
   DFF_X1 \o_buffer_reg[44][13]  (.D(n_132_733), .CK(n_120), .Q(
      \o_buffer[44] [13]), .QN());
   DFF_X1 \o_buffer_reg[44][12]  (.D(n_132_732), .CK(n_120), .Q(
      \o_buffer[44] [12]), .QN());
   DFF_X1 \o_buffer_reg[44][11]  (.D(n_132_731), .CK(n_120), .Q(
      \o_buffer[44] [11]), .QN());
   DFF_X1 \o_buffer_reg[44][10]  (.D(n_132_730), .CK(n_120), .Q(
      \o_buffer[44] [10]), .QN());
   DFF_X1 \o_buffer_reg[44][9]  (.D(n_132_729), .CK(n_120), .Q(\o_buffer[44] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][8]  (.D(n_132_728), .CK(n_120), .Q(\o_buffer[44] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][7]  (.D(n_132_727), .CK(n_120), .Q(\o_buffer[44] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][6]  (.D(n_132_726), .CK(n_120), .Q(\o_buffer[44] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][5]  (.D(n_132_725), .CK(n_120), .Q(\o_buffer[44] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][4]  (.D(n_132_724), .CK(n_120), .Q(\o_buffer[44] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][3]  (.D(n_132_723), .CK(n_120), .Q(\o_buffer[44] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][2]  (.D(n_132_722), .CK(n_120), .Q(\o_buffer[44] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][1]  (.D(n_132_721), .CK(n_120), .Q(\o_buffer[44] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[44][0]  (.D(n_132_720), .CK(n_120), .Q(\o_buffer[44] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][15]  (.D(n_132_719), .CK(n_120), .Q(
      \o_buffer[43] [15]), .QN());
   DFF_X1 \o_buffer_reg[43][14]  (.D(n_132_718), .CK(n_120), .Q(
      \o_buffer[43] [14]), .QN());
   DFF_X1 \o_buffer_reg[43][13]  (.D(n_132_717), .CK(n_120), .Q(
      \o_buffer[43] [13]), .QN());
   DFF_X1 \o_buffer_reg[43][12]  (.D(n_132_716), .CK(n_120), .Q(
      \o_buffer[43] [12]), .QN());
   DFF_X1 \o_buffer_reg[43][11]  (.D(n_132_715), .CK(n_120), .Q(
      \o_buffer[43] [11]), .QN());
   DFF_X1 \o_buffer_reg[43][10]  (.D(n_132_714), .CK(n_120), .Q(
      \o_buffer[43] [10]), .QN());
   DFF_X1 \o_buffer_reg[43][9]  (.D(n_132_713), .CK(n_120), .Q(\o_buffer[43] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][8]  (.D(n_132_712), .CK(n_120), .Q(\o_buffer[43] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][7]  (.D(n_132_711), .CK(n_120), .Q(\o_buffer[43] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][6]  (.D(n_132_710), .CK(n_120), .Q(\o_buffer[43] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][5]  (.D(n_132_709), .CK(n_120), .Q(\o_buffer[43] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][4]  (.D(n_132_708), .CK(n_120), .Q(\o_buffer[43] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][3]  (.D(n_132_707), .CK(n_120), .Q(\o_buffer[43] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][2]  (.D(n_132_706), .CK(n_120), .Q(\o_buffer[43] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][1]  (.D(n_132_705), .CK(n_120), .Q(\o_buffer[43] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[43][0]  (.D(n_132_704), .CK(n_120), .Q(\o_buffer[43] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][15]  (.D(n_132_703), .CK(n_120), .Q(
      \o_buffer[42] [15]), .QN());
   DFF_X1 \o_buffer_reg[42][14]  (.D(n_132_702), .CK(n_120), .Q(
      \o_buffer[42] [14]), .QN());
   DFF_X1 \o_buffer_reg[42][13]  (.D(n_132_701), .CK(n_120), .Q(
      \o_buffer[42] [13]), .QN());
   DFF_X1 \o_buffer_reg[42][12]  (.D(n_132_700), .CK(n_120), .Q(
      \o_buffer[42] [12]), .QN());
   DFF_X1 \o_buffer_reg[42][11]  (.D(n_132_699), .CK(n_120), .Q(
      \o_buffer[42] [11]), .QN());
   DFF_X1 \o_buffer_reg[42][10]  (.D(n_132_698), .CK(n_120), .Q(
      \o_buffer[42] [10]), .QN());
   DFF_X1 \o_buffer_reg[42][9]  (.D(n_132_697), .CK(n_120), .Q(\o_buffer[42] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][8]  (.D(n_132_696), .CK(n_120), .Q(\o_buffer[42] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][7]  (.D(n_132_695), .CK(n_120), .Q(\o_buffer[42] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][6]  (.D(n_132_694), .CK(n_120), .Q(\o_buffer[42] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][5]  (.D(n_132_693), .CK(n_120), .Q(\o_buffer[42] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][4]  (.D(n_132_692), .CK(n_120), .Q(\o_buffer[42] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][3]  (.D(n_132_691), .CK(n_120), .Q(\o_buffer[42] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][2]  (.D(n_132_690), .CK(n_120), .Q(\o_buffer[42] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][1]  (.D(n_132_689), .CK(n_120), .Q(\o_buffer[42] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[42][0]  (.D(n_132_688), .CK(n_120), .Q(\o_buffer[42] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][15]  (.D(n_132_687), .CK(n_120), .Q(
      \o_buffer[41] [15]), .QN());
   DFF_X1 \o_buffer_reg[41][14]  (.D(n_132_686), .CK(n_120), .Q(
      \o_buffer[41] [14]), .QN());
   DFF_X1 \o_buffer_reg[41][13]  (.D(n_132_685), .CK(n_120), .Q(
      \o_buffer[41] [13]), .QN());
   DFF_X1 \o_buffer_reg[41][12]  (.D(n_132_684), .CK(n_120), .Q(
      \o_buffer[41] [12]), .QN());
   DFF_X1 \o_buffer_reg[41][11]  (.D(n_132_683), .CK(n_120), .Q(
      \o_buffer[41] [11]), .QN());
   DFF_X1 \o_buffer_reg[41][10]  (.D(n_132_682), .CK(n_120), .Q(
      \o_buffer[41] [10]), .QN());
   DFF_X1 \o_buffer_reg[41][9]  (.D(n_132_681), .CK(n_120), .Q(\o_buffer[41] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][8]  (.D(n_132_680), .CK(n_120), .Q(\o_buffer[41] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][7]  (.D(n_132_679), .CK(n_120), .Q(\o_buffer[41] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][6]  (.D(n_132_678), .CK(n_120), .Q(\o_buffer[41] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][5]  (.D(n_132_677), .CK(n_120), .Q(\o_buffer[41] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][4]  (.D(n_132_676), .CK(n_120), .Q(\o_buffer[41] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][3]  (.D(n_132_675), .CK(n_120), .Q(\o_buffer[41] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][2]  (.D(n_132_674), .CK(n_120), .Q(\o_buffer[41] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][1]  (.D(n_132_673), .CK(n_120), .Q(\o_buffer[41] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[41][0]  (.D(n_132_672), .CK(n_120), .Q(\o_buffer[41] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][15]  (.D(n_132_671), .CK(n_120), .Q(
      \o_buffer[40] [15]), .QN());
   DFF_X1 \o_buffer_reg[40][14]  (.D(n_132_670), .CK(n_120), .Q(
      \o_buffer[40] [14]), .QN());
   DFF_X1 \o_buffer_reg[40][13]  (.D(n_132_669), .CK(n_120), .Q(
      \o_buffer[40] [13]), .QN());
   DFF_X1 \o_buffer_reg[40][12]  (.D(n_132_668), .CK(n_120), .Q(
      \o_buffer[40] [12]), .QN());
   DFF_X1 \o_buffer_reg[40][11]  (.D(n_132_667), .CK(n_120), .Q(
      \o_buffer[40] [11]), .QN());
   DFF_X1 \o_buffer_reg[40][10]  (.D(n_132_666), .CK(n_120), .Q(
      \o_buffer[40] [10]), .QN());
   DFF_X1 \o_buffer_reg[40][9]  (.D(n_132_665), .CK(n_120), .Q(\o_buffer[40] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][8]  (.D(n_132_664), .CK(n_120), .Q(\o_buffer[40] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][7]  (.D(n_132_663), .CK(n_120), .Q(\o_buffer[40] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][6]  (.D(n_132_662), .CK(n_120), .Q(\o_buffer[40] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][5]  (.D(n_132_661), .CK(n_120), .Q(\o_buffer[40] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][4]  (.D(n_132_660), .CK(n_120), .Q(\o_buffer[40] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][3]  (.D(n_132_659), .CK(n_120), .Q(\o_buffer[40] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][2]  (.D(n_132_658), .CK(n_120), .Q(\o_buffer[40] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][1]  (.D(n_132_657), .CK(n_120), .Q(\o_buffer[40] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[40][0]  (.D(n_132_656), .CK(n_120), .Q(\o_buffer[40] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][15]  (.D(n_132_655), .CK(n_120), .Q(
      \o_buffer[39] [15]), .QN());
   DFF_X1 \o_buffer_reg[39][14]  (.D(n_132_654), .CK(n_120), .Q(
      \o_buffer[39] [14]), .QN());
   DFF_X1 \o_buffer_reg[39][13]  (.D(n_132_653), .CK(n_120), .Q(
      \o_buffer[39] [13]), .QN());
   DFF_X1 \o_buffer_reg[39][12]  (.D(n_132_652), .CK(n_120), .Q(
      \o_buffer[39] [12]), .QN());
   DFF_X1 \o_buffer_reg[39][11]  (.D(n_132_651), .CK(n_120), .Q(
      \o_buffer[39] [11]), .QN());
   DFF_X1 \o_buffer_reg[39][10]  (.D(n_132_650), .CK(n_120), .Q(
      \o_buffer[39] [10]), .QN());
   DFF_X1 \o_buffer_reg[39][9]  (.D(n_132_649), .CK(n_120), .Q(\o_buffer[39] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][8]  (.D(n_132_648), .CK(n_120), .Q(\o_buffer[39] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][7]  (.D(n_132_647), .CK(n_120), .Q(\o_buffer[39] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][6]  (.D(n_132_646), .CK(n_120), .Q(\o_buffer[39] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][5]  (.D(n_132_645), .CK(n_120), .Q(\o_buffer[39] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][4]  (.D(n_132_644), .CK(n_120), .Q(\o_buffer[39] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][3]  (.D(n_132_643), .CK(n_120), .Q(\o_buffer[39] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][2]  (.D(n_132_642), .CK(n_120), .Q(\o_buffer[39] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][1]  (.D(n_132_641), .CK(n_120), .Q(\o_buffer[39] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[39][0]  (.D(n_132_640), .CK(n_120), .Q(\o_buffer[39] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][15]  (.D(n_132_639), .CK(n_120), .Q(
      \o_buffer[38] [15]), .QN());
   DFF_X1 \o_buffer_reg[38][14]  (.D(n_132_638), .CK(n_120), .Q(
      \o_buffer[38] [14]), .QN());
   DFF_X1 \o_buffer_reg[38][13]  (.D(n_132_637), .CK(n_120), .Q(
      \o_buffer[38] [13]), .QN());
   DFF_X1 \o_buffer_reg[38][12]  (.D(n_132_636), .CK(n_120), .Q(
      \o_buffer[38] [12]), .QN());
   DFF_X1 \o_buffer_reg[38][11]  (.D(n_132_635), .CK(n_120), .Q(
      \o_buffer[38] [11]), .QN());
   DFF_X1 \o_buffer_reg[38][10]  (.D(n_132_634), .CK(n_120), .Q(
      \o_buffer[38] [10]), .QN());
   DFF_X1 \o_buffer_reg[38][9]  (.D(n_132_633), .CK(n_120), .Q(\o_buffer[38] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][8]  (.D(n_132_632), .CK(n_120), .Q(\o_buffer[38] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][7]  (.D(n_132_631), .CK(n_120), .Q(\o_buffer[38] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][6]  (.D(n_132_630), .CK(n_120), .Q(\o_buffer[38] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][5]  (.D(n_132_629), .CK(n_120), .Q(\o_buffer[38] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][4]  (.D(n_132_628), .CK(n_120), .Q(\o_buffer[38] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][3]  (.D(n_132_627), .CK(n_120), .Q(\o_buffer[38] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][2]  (.D(n_132_626), .CK(n_120), .Q(\o_buffer[38] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][1]  (.D(n_132_625), .CK(n_120), .Q(\o_buffer[38] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[38][0]  (.D(n_132_624), .CK(n_120), .Q(\o_buffer[38] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][15]  (.D(n_132_623), .CK(n_120), .Q(
      \o_buffer[37] [15]), .QN());
   DFF_X1 \o_buffer_reg[37][14]  (.D(n_132_622), .CK(n_120), .Q(
      \o_buffer[37] [14]), .QN());
   DFF_X1 \o_buffer_reg[37][13]  (.D(n_132_621), .CK(n_120), .Q(
      \o_buffer[37] [13]), .QN());
   DFF_X1 \o_buffer_reg[37][12]  (.D(n_132_620), .CK(n_120), .Q(
      \o_buffer[37] [12]), .QN());
   DFF_X1 \o_buffer_reg[37][11]  (.D(n_132_619), .CK(n_120), .Q(
      \o_buffer[37] [11]), .QN());
   DFF_X1 \o_buffer_reg[37][10]  (.D(n_132_618), .CK(n_120), .Q(
      \o_buffer[37] [10]), .QN());
   DFF_X1 \o_buffer_reg[37][9]  (.D(n_132_617), .CK(n_120), .Q(\o_buffer[37] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][8]  (.D(n_132_616), .CK(n_120), .Q(\o_buffer[37] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][7]  (.D(n_132_615), .CK(n_120), .Q(\o_buffer[37] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][6]  (.D(n_132_614), .CK(n_120), .Q(\o_buffer[37] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][5]  (.D(n_132_613), .CK(n_120), .Q(\o_buffer[37] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][4]  (.D(n_132_612), .CK(n_120), .Q(\o_buffer[37] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][3]  (.D(n_132_611), .CK(n_120), .Q(\o_buffer[37] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][2]  (.D(n_132_610), .CK(n_120), .Q(\o_buffer[37] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][1]  (.D(n_132_609), .CK(n_120), .Q(\o_buffer[37] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[37][0]  (.D(n_132_608), .CK(n_120), .Q(\o_buffer[37] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][15]  (.D(n_132_607), .CK(n_120), .Q(
      \o_buffer[36] [15]), .QN());
   DFF_X1 \o_buffer_reg[36][14]  (.D(n_132_606), .CK(n_120), .Q(
      \o_buffer[36] [14]), .QN());
   DFF_X1 \o_buffer_reg[36][13]  (.D(n_132_605), .CK(n_120), .Q(
      \o_buffer[36] [13]), .QN());
   DFF_X1 \o_buffer_reg[36][12]  (.D(n_132_604), .CK(n_120), .Q(
      \o_buffer[36] [12]), .QN());
   DFF_X1 \o_buffer_reg[36][11]  (.D(n_132_603), .CK(n_120), .Q(
      \o_buffer[36] [11]), .QN());
   DFF_X1 \o_buffer_reg[36][10]  (.D(n_132_602), .CK(n_120), .Q(
      \o_buffer[36] [10]), .QN());
   DFF_X1 \o_buffer_reg[36][9]  (.D(n_132_601), .CK(n_120), .Q(\o_buffer[36] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][8]  (.D(n_132_600), .CK(n_120), .Q(\o_buffer[36] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][7]  (.D(n_132_599), .CK(n_120), .Q(\o_buffer[36] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][6]  (.D(n_132_598), .CK(n_120), .Q(\o_buffer[36] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][5]  (.D(n_132_597), .CK(n_120), .Q(\o_buffer[36] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][4]  (.D(n_132_596), .CK(n_120), .Q(\o_buffer[36] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][3]  (.D(n_132_595), .CK(n_120), .Q(\o_buffer[36] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][2]  (.D(n_132_594), .CK(n_120), .Q(\o_buffer[36] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][1]  (.D(n_132_593), .CK(n_120), .Q(\o_buffer[36] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[36][0]  (.D(n_132_592), .CK(n_120), .Q(\o_buffer[36] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][15]  (.D(n_132_591), .CK(n_120), .Q(
      \o_buffer[35] [15]), .QN());
   DFF_X1 \o_buffer_reg[35][14]  (.D(n_132_590), .CK(n_120), .Q(
      \o_buffer[35] [14]), .QN());
   DFF_X1 \o_buffer_reg[35][13]  (.D(n_132_589), .CK(n_120), .Q(
      \o_buffer[35] [13]), .QN());
   DFF_X1 \o_buffer_reg[35][12]  (.D(n_132_588), .CK(n_120), .Q(
      \o_buffer[35] [12]), .QN());
   DFF_X1 \o_buffer_reg[35][11]  (.D(n_132_587), .CK(n_120), .Q(
      \o_buffer[35] [11]), .QN());
   DFF_X1 \o_buffer_reg[35][10]  (.D(n_132_586), .CK(n_120), .Q(
      \o_buffer[35] [10]), .QN());
   DFF_X1 \o_buffer_reg[35][9]  (.D(n_132_585), .CK(n_120), .Q(\o_buffer[35] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][8]  (.D(n_132_584), .CK(n_120), .Q(\o_buffer[35] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][7]  (.D(n_132_583), .CK(n_120), .Q(\o_buffer[35] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][6]  (.D(n_132_582), .CK(n_120), .Q(\o_buffer[35] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][5]  (.D(n_132_581), .CK(n_120), .Q(\o_buffer[35] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][4]  (.D(n_132_580), .CK(n_120), .Q(\o_buffer[35] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][3]  (.D(n_132_579), .CK(n_120), .Q(\o_buffer[35] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][2]  (.D(n_132_578), .CK(n_120), .Q(\o_buffer[35] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][1]  (.D(n_132_577), .CK(n_120), .Q(\o_buffer[35] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[35][0]  (.D(n_132_576), .CK(n_120), .Q(\o_buffer[35] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][15]  (.D(n_132_575), .CK(n_120), .Q(
      \o_buffer[34] [15]), .QN());
   DFF_X1 \o_buffer_reg[34][14]  (.D(n_132_574), .CK(n_120), .Q(
      \o_buffer[34] [14]), .QN());
   DFF_X1 \o_buffer_reg[34][13]  (.D(n_132_573), .CK(n_120), .Q(
      \o_buffer[34] [13]), .QN());
   DFF_X1 \o_buffer_reg[34][12]  (.D(n_132_572), .CK(n_120), .Q(
      \o_buffer[34] [12]), .QN());
   DFF_X1 \o_buffer_reg[34][11]  (.D(n_132_571), .CK(n_120), .Q(
      \o_buffer[34] [11]), .QN());
   DFF_X1 \o_buffer_reg[34][10]  (.D(n_132_570), .CK(n_120), .Q(
      \o_buffer[34] [10]), .QN());
   DFF_X1 \o_buffer_reg[34][9]  (.D(n_132_569), .CK(n_120), .Q(\o_buffer[34] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][8]  (.D(n_132_568), .CK(n_120), .Q(\o_buffer[34] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][7]  (.D(n_132_567), .CK(n_120), .Q(\o_buffer[34] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][6]  (.D(n_132_566), .CK(n_120), .Q(\o_buffer[34] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][5]  (.D(n_132_565), .CK(n_120), .Q(\o_buffer[34] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][4]  (.D(n_132_564), .CK(n_120), .Q(\o_buffer[34] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][3]  (.D(n_132_563), .CK(n_120), .Q(\o_buffer[34] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][2]  (.D(n_132_562), .CK(n_120), .Q(\o_buffer[34] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][1]  (.D(n_132_561), .CK(n_120), .Q(\o_buffer[34] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[34][0]  (.D(n_132_560), .CK(n_120), .Q(\o_buffer[34] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][15]  (.D(n_132_559), .CK(n_120), .Q(
      \o_buffer[33] [15]), .QN());
   DFF_X1 \o_buffer_reg[33][14]  (.D(n_132_558), .CK(n_120), .Q(
      \o_buffer[33] [14]), .QN());
   DFF_X1 \o_buffer_reg[33][13]  (.D(n_132_557), .CK(n_120), .Q(
      \o_buffer[33] [13]), .QN());
   DFF_X1 \o_buffer_reg[33][12]  (.D(n_132_556), .CK(n_120), .Q(
      \o_buffer[33] [12]), .QN());
   DFF_X1 \o_buffer_reg[33][11]  (.D(n_132_555), .CK(n_120), .Q(
      \o_buffer[33] [11]), .QN());
   DFF_X1 \o_buffer_reg[33][10]  (.D(n_132_554), .CK(n_120), .Q(
      \o_buffer[33] [10]), .QN());
   DFF_X1 \o_buffer_reg[33][9]  (.D(n_132_553), .CK(n_120), .Q(\o_buffer[33] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][8]  (.D(n_132_552), .CK(n_120), .Q(\o_buffer[33] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][7]  (.D(n_132_551), .CK(n_120), .Q(\o_buffer[33] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][6]  (.D(n_132_550), .CK(n_120), .Q(\o_buffer[33] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][5]  (.D(n_132_549), .CK(n_120), .Q(\o_buffer[33] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][4]  (.D(n_132_548), .CK(n_120), .Q(\o_buffer[33] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][3]  (.D(n_132_547), .CK(n_120), .Q(\o_buffer[33] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][2]  (.D(n_132_546), .CK(n_120), .Q(\o_buffer[33] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][1]  (.D(n_132_545), .CK(n_120), .Q(\o_buffer[33] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[33][0]  (.D(n_132_544), .CK(n_120), .Q(\o_buffer[33] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][15]  (.D(n_132_543), .CK(n_120), .Q(
      \o_buffer[32] [15]), .QN());
   DFF_X1 \o_buffer_reg[32][14]  (.D(n_132_542), .CK(n_120), .Q(
      \o_buffer[32] [14]), .QN());
   DFF_X1 \o_buffer_reg[32][13]  (.D(n_132_541), .CK(n_120), .Q(
      \o_buffer[32] [13]), .QN());
   DFF_X1 \o_buffer_reg[32][12]  (.D(n_132_540), .CK(n_120), .Q(
      \o_buffer[32] [12]), .QN());
   DFF_X1 \o_buffer_reg[32][11]  (.D(n_132_539), .CK(n_120), .Q(
      \o_buffer[32] [11]), .QN());
   DFF_X1 \o_buffer_reg[32][10]  (.D(n_132_538), .CK(n_120), .Q(
      \o_buffer[32] [10]), .QN());
   DFF_X1 \o_buffer_reg[32][9]  (.D(n_132_537), .CK(n_120), .Q(\o_buffer[32] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][8]  (.D(n_132_536), .CK(n_120), .Q(\o_buffer[32] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][7]  (.D(n_132_535), .CK(n_120), .Q(\o_buffer[32] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][6]  (.D(n_132_534), .CK(n_120), .Q(\o_buffer[32] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][5]  (.D(n_132_533), .CK(n_120), .Q(\o_buffer[32] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][4]  (.D(n_132_532), .CK(n_120), .Q(\o_buffer[32] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][3]  (.D(n_132_531), .CK(n_120), .Q(\o_buffer[32] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][2]  (.D(n_132_530), .CK(n_120), .Q(\o_buffer[32] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][1]  (.D(n_132_529), .CK(n_120), .Q(\o_buffer[32] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[32][0]  (.D(n_132_528), .CK(n_120), .Q(\o_buffer[32] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][15]  (.D(n_132_527), .CK(n_120), .Q(
      \o_buffer[31] [15]), .QN());
   DFF_X1 \o_buffer_reg[31][14]  (.D(n_132_526), .CK(n_120), .Q(
      \o_buffer[31] [14]), .QN());
   DFF_X1 \o_buffer_reg[31][13]  (.D(n_132_525), .CK(n_120), .Q(
      \o_buffer[31] [13]), .QN());
   DFF_X1 \o_buffer_reg[31][12]  (.D(n_132_524), .CK(n_120), .Q(
      \o_buffer[31] [12]), .QN());
   DFF_X1 \o_buffer_reg[31][11]  (.D(n_132_523), .CK(n_120), .Q(
      \o_buffer[31] [11]), .QN());
   DFF_X1 \o_buffer_reg[31][10]  (.D(n_132_522), .CK(n_120), .Q(
      \o_buffer[31] [10]), .QN());
   DFF_X1 \o_buffer_reg[31][9]  (.D(n_132_521), .CK(n_120), .Q(\o_buffer[31] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][8]  (.D(n_132_520), .CK(n_120), .Q(\o_buffer[31] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][7]  (.D(n_132_519), .CK(n_120), .Q(\o_buffer[31] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][6]  (.D(n_132_518), .CK(n_120), .Q(\o_buffer[31] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][5]  (.D(n_132_517), .CK(n_120), .Q(\o_buffer[31] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][4]  (.D(n_132_516), .CK(n_120), .Q(\o_buffer[31] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][3]  (.D(n_132_515), .CK(n_120), .Q(\o_buffer[31] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][2]  (.D(n_132_514), .CK(n_120), .Q(\o_buffer[31] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][1]  (.D(n_132_513), .CK(n_120), .Q(\o_buffer[31] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[31][0]  (.D(n_132_512), .CK(n_120), .Q(\o_buffer[31] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][15]  (.D(n_132_511), .CK(n_120), .Q(
      \o_buffer[30] [15]), .QN());
   DFF_X1 \o_buffer_reg[30][14]  (.D(n_132_510), .CK(n_120), .Q(
      \o_buffer[30] [14]), .QN());
   DFF_X1 \o_buffer_reg[30][13]  (.D(n_132_509), .CK(n_120), .Q(
      \o_buffer[30] [13]), .QN());
   DFF_X1 \o_buffer_reg[30][12]  (.D(n_132_508), .CK(n_120), .Q(
      \o_buffer[30] [12]), .QN());
   DFF_X1 \o_buffer_reg[30][11]  (.D(n_132_507), .CK(n_120), .Q(
      \o_buffer[30] [11]), .QN());
   DFF_X1 \o_buffer_reg[30][10]  (.D(n_132_506), .CK(n_120), .Q(
      \o_buffer[30] [10]), .QN());
   DFF_X1 \o_buffer_reg[30][9]  (.D(n_132_505), .CK(n_120), .Q(\o_buffer[30] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][8]  (.D(n_132_504), .CK(n_120), .Q(\o_buffer[30] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][7]  (.D(n_132_503), .CK(n_120), .Q(\o_buffer[30] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][6]  (.D(n_132_502), .CK(n_120), .Q(\o_buffer[30] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][5]  (.D(n_132_501), .CK(n_120), .Q(\o_buffer[30] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][4]  (.D(n_132_500), .CK(n_120), .Q(\o_buffer[30] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][3]  (.D(n_132_499), .CK(n_120), .Q(\o_buffer[30] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][2]  (.D(n_132_498), .CK(n_120), .Q(\o_buffer[30] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][1]  (.D(n_132_497), .CK(n_120), .Q(\o_buffer[30] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[30][0]  (.D(n_132_496), .CK(n_120), .Q(\o_buffer[30] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][15]  (.D(n_132_495), .CK(n_120), .Q(
      \o_buffer[29] [15]), .QN());
   DFF_X1 \o_buffer_reg[29][14]  (.D(n_132_494), .CK(n_120), .Q(
      \o_buffer[29] [14]), .QN());
   DFF_X1 \o_buffer_reg[29][13]  (.D(n_132_493), .CK(n_120), .Q(
      \o_buffer[29] [13]), .QN());
   DFF_X1 \o_buffer_reg[29][12]  (.D(n_132_492), .CK(n_120), .Q(
      \o_buffer[29] [12]), .QN());
   DFF_X1 \o_buffer_reg[29][11]  (.D(n_132_491), .CK(n_120), .Q(
      \o_buffer[29] [11]), .QN());
   DFF_X1 \o_buffer_reg[29][10]  (.D(n_132_490), .CK(n_120), .Q(
      \o_buffer[29] [10]), .QN());
   DFF_X1 \o_buffer_reg[29][9]  (.D(n_132_489), .CK(n_120), .Q(\o_buffer[29] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][8]  (.D(n_132_488), .CK(n_120), .Q(\o_buffer[29] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][7]  (.D(n_132_487), .CK(n_120), .Q(\o_buffer[29] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][6]  (.D(n_132_486), .CK(n_120), .Q(\o_buffer[29] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][5]  (.D(n_132_485), .CK(n_120), .Q(\o_buffer[29] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][4]  (.D(n_132_484), .CK(n_120), .Q(\o_buffer[29] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][3]  (.D(n_132_483), .CK(n_120), .Q(\o_buffer[29] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][2]  (.D(n_132_482), .CK(n_120), .Q(\o_buffer[29] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][1]  (.D(n_132_481), .CK(n_120), .Q(\o_buffer[29] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[29][0]  (.D(n_132_480), .CK(n_120), .Q(\o_buffer[29] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][15]  (.D(n_132_479), .CK(n_120), .Q(
      \o_buffer[28] [15]), .QN());
   DFF_X1 \o_buffer_reg[28][14]  (.D(n_132_478), .CK(n_120), .Q(
      \o_buffer[28] [14]), .QN());
   DFF_X1 \o_buffer_reg[28][13]  (.D(n_132_477), .CK(n_120), .Q(
      \o_buffer[28] [13]), .QN());
   DFF_X1 \o_buffer_reg[28][12]  (.D(n_132_476), .CK(n_120), .Q(
      \o_buffer[28] [12]), .QN());
   DFF_X1 \o_buffer_reg[28][11]  (.D(n_132_475), .CK(n_120), .Q(
      \o_buffer[28] [11]), .QN());
   DFF_X1 \o_buffer_reg[28][10]  (.D(n_132_474), .CK(n_120), .Q(
      \o_buffer[28] [10]), .QN());
   DFF_X1 \o_buffer_reg[28][9]  (.D(n_132_473), .CK(n_120), .Q(\o_buffer[28] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][8]  (.D(n_132_472), .CK(n_120), .Q(\o_buffer[28] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][7]  (.D(n_132_471), .CK(n_120), .Q(\o_buffer[28] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][6]  (.D(n_132_470), .CK(n_120), .Q(\o_buffer[28] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][5]  (.D(n_132_469), .CK(n_120), .Q(\o_buffer[28] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][4]  (.D(n_132_468), .CK(n_120), .Q(\o_buffer[28] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][3]  (.D(n_132_467), .CK(n_120), .Q(\o_buffer[28] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][2]  (.D(n_132_466), .CK(n_120), .Q(\o_buffer[28] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][1]  (.D(n_132_465), .CK(n_120), .Q(\o_buffer[28] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[28][0]  (.D(n_132_464), .CK(n_120), .Q(\o_buffer[28] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][15]  (.D(n_132_463), .CK(n_120), .Q(
      \o_buffer[27] [15]), .QN());
   DFF_X1 \o_buffer_reg[27][14]  (.D(n_132_462), .CK(n_120), .Q(
      \o_buffer[27] [14]), .QN());
   DFF_X1 \o_buffer_reg[27][13]  (.D(n_132_461), .CK(n_120), .Q(
      \o_buffer[27] [13]), .QN());
   DFF_X1 \o_buffer_reg[27][12]  (.D(n_132_460), .CK(n_120), .Q(
      \o_buffer[27] [12]), .QN());
   DFF_X1 \o_buffer_reg[27][11]  (.D(n_132_459), .CK(n_120), .Q(
      \o_buffer[27] [11]), .QN());
   DFF_X1 \o_buffer_reg[27][10]  (.D(n_132_458), .CK(n_120), .Q(
      \o_buffer[27] [10]), .QN());
   DFF_X1 \o_buffer_reg[27][9]  (.D(n_132_457), .CK(n_120), .Q(\o_buffer[27] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][8]  (.D(n_132_456), .CK(n_120), .Q(\o_buffer[27] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][7]  (.D(n_132_455), .CK(n_120), .Q(\o_buffer[27] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][6]  (.D(n_132_454), .CK(n_120), .Q(\o_buffer[27] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][5]  (.D(n_132_453), .CK(n_120), .Q(\o_buffer[27] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][4]  (.D(n_132_452), .CK(n_120), .Q(\o_buffer[27] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][3]  (.D(n_132_451), .CK(n_120), .Q(\o_buffer[27] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][2]  (.D(n_132_450), .CK(n_120), .Q(\o_buffer[27] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][1]  (.D(n_132_449), .CK(n_120), .Q(\o_buffer[27] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[27][0]  (.D(n_132_448), .CK(n_120), .Q(\o_buffer[27] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][15]  (.D(n_132_447), .CK(n_120), .Q(
      \o_buffer[26] [15]), .QN());
   DFF_X1 \o_buffer_reg[26][14]  (.D(n_132_446), .CK(n_120), .Q(
      \o_buffer[26] [14]), .QN());
   DFF_X1 \o_buffer_reg[26][13]  (.D(n_132_445), .CK(n_120), .Q(
      \o_buffer[26] [13]), .QN());
   DFF_X1 \o_buffer_reg[26][12]  (.D(n_132_444), .CK(n_120), .Q(
      \o_buffer[26] [12]), .QN());
   DFF_X1 \o_buffer_reg[26][11]  (.D(n_132_443), .CK(n_120), .Q(
      \o_buffer[26] [11]), .QN());
   DFF_X1 \o_buffer_reg[26][10]  (.D(n_132_442), .CK(n_120), .Q(
      \o_buffer[26] [10]), .QN());
   DFF_X1 \o_buffer_reg[26][9]  (.D(n_132_441), .CK(n_120), .Q(\o_buffer[26] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][8]  (.D(n_132_440), .CK(n_120), .Q(\o_buffer[26] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][7]  (.D(n_132_439), .CK(n_120), .Q(\o_buffer[26] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][6]  (.D(n_132_438), .CK(n_120), .Q(\o_buffer[26] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][5]  (.D(n_132_437), .CK(n_120), .Q(\o_buffer[26] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][4]  (.D(n_132_436), .CK(n_120), .Q(\o_buffer[26] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][3]  (.D(n_132_435), .CK(n_120), .Q(\o_buffer[26] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][2]  (.D(n_132_434), .CK(n_120), .Q(\o_buffer[26] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][1]  (.D(n_132_433), .CK(n_120), .Q(\o_buffer[26] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[26][0]  (.D(n_132_432), .CK(n_120), .Q(\o_buffer[26] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][15]  (.D(n_132_431), .CK(n_120), .Q(
      \o_buffer[25] [15]), .QN());
   DFF_X1 \o_buffer_reg[25][14]  (.D(n_132_430), .CK(n_120), .Q(
      \o_buffer[25] [14]), .QN());
   DFF_X1 \o_buffer_reg[25][13]  (.D(n_132_429), .CK(n_120), .Q(
      \o_buffer[25] [13]), .QN());
   DFF_X1 \o_buffer_reg[25][12]  (.D(n_132_428), .CK(n_120), .Q(
      \o_buffer[25] [12]), .QN());
   DFF_X1 \o_buffer_reg[25][11]  (.D(n_132_427), .CK(n_120), .Q(
      \o_buffer[25] [11]), .QN());
   DFF_X1 \o_buffer_reg[25][10]  (.D(n_132_426), .CK(n_120), .Q(
      \o_buffer[25] [10]), .QN());
   DFF_X1 \o_buffer_reg[25][9]  (.D(n_132_425), .CK(n_120), .Q(\o_buffer[25] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][8]  (.D(n_132_424), .CK(n_120), .Q(\o_buffer[25] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][7]  (.D(n_132_423), .CK(n_120), .Q(\o_buffer[25] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][6]  (.D(n_132_422), .CK(n_120), .Q(\o_buffer[25] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][5]  (.D(n_132_421), .CK(n_120), .Q(\o_buffer[25] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][4]  (.D(n_132_420), .CK(n_120), .Q(\o_buffer[25] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][3]  (.D(n_132_419), .CK(n_120), .Q(\o_buffer[25] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][2]  (.D(n_132_418), .CK(n_120), .Q(\o_buffer[25] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][1]  (.D(n_132_417), .CK(n_120), .Q(\o_buffer[25] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[25][0]  (.D(n_132_416), .CK(n_120), .Q(\o_buffer[25] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][15]  (.D(n_132_415), .CK(n_120), .Q(
      \o_buffer[24] [15]), .QN());
   DFF_X1 \o_buffer_reg[24][14]  (.D(n_132_414), .CK(n_120), .Q(
      \o_buffer[24] [14]), .QN());
   DFF_X1 \o_buffer_reg[24][13]  (.D(n_132_413), .CK(n_120), .Q(
      \o_buffer[24] [13]), .QN());
   DFF_X1 \o_buffer_reg[24][12]  (.D(n_132_412), .CK(n_120), .Q(
      \o_buffer[24] [12]), .QN());
   DFF_X1 \o_buffer_reg[24][11]  (.D(n_132_411), .CK(n_120), .Q(
      \o_buffer[24] [11]), .QN());
   DFF_X1 \o_buffer_reg[24][10]  (.D(n_132_410), .CK(n_120), .Q(
      \o_buffer[24] [10]), .QN());
   DFF_X1 \o_buffer_reg[24][9]  (.D(n_132_409), .CK(n_120), .Q(\o_buffer[24] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][8]  (.D(n_132_408), .CK(n_120), .Q(\o_buffer[24] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][7]  (.D(n_132_407), .CK(n_120), .Q(\o_buffer[24] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][6]  (.D(n_132_406), .CK(n_120), .Q(\o_buffer[24] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][5]  (.D(n_132_405), .CK(n_120), .Q(\o_buffer[24] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][4]  (.D(n_132_404), .CK(n_120), .Q(\o_buffer[24] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][3]  (.D(n_132_403), .CK(n_120), .Q(\o_buffer[24] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][2]  (.D(n_132_402), .CK(n_120), .Q(\o_buffer[24] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][1]  (.D(n_132_401), .CK(n_120), .Q(\o_buffer[24] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[24][0]  (.D(n_132_400), .CK(n_120), .Q(\o_buffer[24] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][15]  (.D(n_132_399), .CK(n_120), .Q(
      \o_buffer[23] [15]), .QN());
   DFF_X1 \o_buffer_reg[23][14]  (.D(n_132_398), .CK(n_120), .Q(
      \o_buffer[23] [14]), .QN());
   DFF_X1 \o_buffer_reg[23][13]  (.D(n_132_397), .CK(n_120), .Q(
      \o_buffer[23] [13]), .QN());
   DFF_X1 \o_buffer_reg[23][12]  (.D(n_132_396), .CK(n_120), .Q(
      \o_buffer[23] [12]), .QN());
   DFF_X1 \o_buffer_reg[23][11]  (.D(n_132_395), .CK(n_120), .Q(
      \o_buffer[23] [11]), .QN());
   DFF_X1 \o_buffer_reg[23][10]  (.D(n_132_394), .CK(n_120), .Q(
      \o_buffer[23] [10]), .QN());
   DFF_X1 \o_buffer_reg[23][9]  (.D(n_132_393), .CK(n_120), .Q(\o_buffer[23] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][8]  (.D(n_132_392), .CK(n_120), .Q(\o_buffer[23] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][7]  (.D(n_132_391), .CK(n_120), .Q(\o_buffer[23] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][6]  (.D(n_132_390), .CK(n_120), .Q(\o_buffer[23] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][5]  (.D(n_132_389), .CK(n_120), .Q(\o_buffer[23] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][4]  (.D(n_132_388), .CK(n_120), .Q(\o_buffer[23] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][3]  (.D(n_132_387), .CK(n_120), .Q(\o_buffer[23] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][2]  (.D(n_132_386), .CK(n_120), .Q(\o_buffer[23] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][1]  (.D(n_132_385), .CK(n_120), .Q(\o_buffer[23] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[23][0]  (.D(n_132_384), .CK(n_120), .Q(\o_buffer[23] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][15]  (.D(n_132_383), .CK(n_120), .Q(
      \o_buffer[22] [15]), .QN());
   DFF_X1 \o_buffer_reg[22][14]  (.D(n_132_382), .CK(n_120), .Q(
      \o_buffer[22] [14]), .QN());
   DFF_X1 \o_buffer_reg[22][13]  (.D(n_132_381), .CK(n_120), .Q(
      \o_buffer[22] [13]), .QN());
   DFF_X1 \o_buffer_reg[22][12]  (.D(n_132_380), .CK(n_120), .Q(
      \o_buffer[22] [12]), .QN());
   DFF_X1 \o_buffer_reg[22][11]  (.D(n_132_379), .CK(n_120), .Q(
      \o_buffer[22] [11]), .QN());
   DFF_X1 \o_buffer_reg[22][10]  (.D(n_132_378), .CK(n_120), .Q(
      \o_buffer[22] [10]), .QN());
   DFF_X1 \o_buffer_reg[22][9]  (.D(n_132_377), .CK(n_120), .Q(\o_buffer[22] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][8]  (.D(n_132_376), .CK(n_120), .Q(\o_buffer[22] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][7]  (.D(n_132_375), .CK(n_120), .Q(\o_buffer[22] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][6]  (.D(n_132_374), .CK(n_120), .Q(\o_buffer[22] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][5]  (.D(n_132_373), .CK(n_120), .Q(\o_buffer[22] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][4]  (.D(n_132_372), .CK(n_120), .Q(\o_buffer[22] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][3]  (.D(n_132_371), .CK(n_120), .Q(\o_buffer[22] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][2]  (.D(n_132_370), .CK(n_120), .Q(\o_buffer[22] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][1]  (.D(n_132_369), .CK(n_120), .Q(\o_buffer[22] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[22][0]  (.D(n_132_368), .CK(n_120), .Q(\o_buffer[22] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][15]  (.D(n_132_367), .CK(n_120), .Q(
      \o_buffer[21] [15]), .QN());
   DFF_X1 \o_buffer_reg[21][14]  (.D(n_132_366), .CK(n_120), .Q(
      \o_buffer[21] [14]), .QN());
   DFF_X1 \o_buffer_reg[21][13]  (.D(n_132_365), .CK(n_120), .Q(
      \o_buffer[21] [13]), .QN());
   DFF_X1 \o_buffer_reg[21][12]  (.D(n_132_364), .CK(n_120), .Q(
      \o_buffer[21] [12]), .QN());
   DFF_X1 \o_buffer_reg[21][11]  (.D(n_132_363), .CK(n_120), .Q(
      \o_buffer[21] [11]), .QN());
   DFF_X1 \o_buffer_reg[21][10]  (.D(n_132_362), .CK(n_120), .Q(
      \o_buffer[21] [10]), .QN());
   DFF_X1 \o_buffer_reg[21][9]  (.D(n_132_361), .CK(n_120), .Q(\o_buffer[21] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][8]  (.D(n_132_360), .CK(n_120), .Q(\o_buffer[21] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][7]  (.D(n_132_359), .CK(n_120), .Q(\o_buffer[21] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][6]  (.D(n_132_358), .CK(n_120), .Q(\o_buffer[21] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][5]  (.D(n_132_357), .CK(n_120), .Q(\o_buffer[21] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][4]  (.D(n_132_356), .CK(n_120), .Q(\o_buffer[21] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][3]  (.D(n_132_355), .CK(n_120), .Q(\o_buffer[21] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][2]  (.D(n_132_354), .CK(n_120), .Q(\o_buffer[21] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][1]  (.D(n_132_353), .CK(n_120), .Q(\o_buffer[21] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[21][0]  (.D(n_132_352), .CK(n_120), .Q(\o_buffer[21] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][15]  (.D(n_132_351), .CK(n_120), .Q(
      \o_buffer[20] [15]), .QN());
   DFF_X1 \o_buffer_reg[20][14]  (.D(n_132_350), .CK(n_120), .Q(
      \o_buffer[20] [14]), .QN());
   DFF_X1 \o_buffer_reg[20][13]  (.D(n_132_349), .CK(n_120), .Q(
      \o_buffer[20] [13]), .QN());
   DFF_X1 \o_buffer_reg[20][12]  (.D(n_132_348), .CK(n_120), .Q(
      \o_buffer[20] [12]), .QN());
   DFF_X1 \o_buffer_reg[20][11]  (.D(n_132_347), .CK(n_120), .Q(
      \o_buffer[20] [11]), .QN());
   DFF_X1 \o_buffer_reg[20][10]  (.D(n_132_346), .CK(n_120), .Q(
      \o_buffer[20] [10]), .QN());
   DFF_X1 \o_buffer_reg[20][9]  (.D(n_132_345), .CK(n_120), .Q(\o_buffer[20] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][8]  (.D(n_132_344), .CK(n_120), .Q(\o_buffer[20] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][7]  (.D(n_132_343), .CK(n_120), .Q(\o_buffer[20] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][6]  (.D(n_132_342), .CK(n_120), .Q(\o_buffer[20] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][5]  (.D(n_132_341), .CK(n_120), .Q(\o_buffer[20] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][4]  (.D(n_132_340), .CK(n_120), .Q(\o_buffer[20] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][3]  (.D(n_132_339), .CK(n_120), .Q(\o_buffer[20] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][2]  (.D(n_132_338), .CK(n_120), .Q(\o_buffer[20] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][1]  (.D(n_132_337), .CK(n_120), .Q(\o_buffer[20] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[20][0]  (.D(n_132_336), .CK(n_120), .Q(\o_buffer[20] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][15]  (.D(n_132_335), .CK(n_120), .Q(
      \o_buffer[19] [15]), .QN());
   DFF_X1 \o_buffer_reg[19][14]  (.D(n_132_334), .CK(n_120), .Q(
      \o_buffer[19] [14]), .QN());
   DFF_X1 \o_buffer_reg[19][13]  (.D(n_132_333), .CK(n_120), .Q(
      \o_buffer[19] [13]), .QN());
   DFF_X1 \o_buffer_reg[19][12]  (.D(n_132_332), .CK(n_120), .Q(
      \o_buffer[19] [12]), .QN());
   DFF_X1 \o_buffer_reg[19][11]  (.D(n_132_331), .CK(n_120), .Q(
      \o_buffer[19] [11]), .QN());
   DFF_X1 \o_buffer_reg[19][10]  (.D(n_132_330), .CK(n_120), .Q(
      \o_buffer[19] [10]), .QN());
   DFF_X1 \o_buffer_reg[19][9]  (.D(n_132_329), .CK(n_120), .Q(\o_buffer[19] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][8]  (.D(n_132_328), .CK(n_120), .Q(\o_buffer[19] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][7]  (.D(n_132_327), .CK(n_120), .Q(\o_buffer[19] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][6]  (.D(n_132_326), .CK(n_120), .Q(\o_buffer[19] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][5]  (.D(n_132_325), .CK(n_120), .Q(\o_buffer[19] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][4]  (.D(n_132_324), .CK(n_120), .Q(\o_buffer[19] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][3]  (.D(n_132_323), .CK(n_120), .Q(\o_buffer[19] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][2]  (.D(n_132_322), .CK(n_120), .Q(\o_buffer[19] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][1]  (.D(n_132_321), .CK(n_120), .Q(\o_buffer[19] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[19][0]  (.D(n_132_320), .CK(n_120), .Q(\o_buffer[19] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][15]  (.D(n_132_319), .CK(n_120), .Q(
      \o_buffer[18] [15]), .QN());
   DFF_X1 \o_buffer_reg[18][14]  (.D(n_132_318), .CK(n_120), .Q(
      \o_buffer[18] [14]), .QN());
   DFF_X1 \o_buffer_reg[18][13]  (.D(n_132_317), .CK(n_120), .Q(
      \o_buffer[18] [13]), .QN());
   DFF_X1 \o_buffer_reg[18][12]  (.D(n_132_316), .CK(n_120), .Q(
      \o_buffer[18] [12]), .QN());
   DFF_X1 \o_buffer_reg[18][11]  (.D(n_132_315), .CK(n_120), .Q(
      \o_buffer[18] [11]), .QN());
   DFF_X1 \o_buffer_reg[18][10]  (.D(n_132_314), .CK(n_120), .Q(
      \o_buffer[18] [10]), .QN());
   DFF_X1 \o_buffer_reg[18][9]  (.D(n_132_313), .CK(n_120), .Q(\o_buffer[18] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][8]  (.D(n_132_312), .CK(n_120), .Q(\o_buffer[18] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][7]  (.D(n_132_311), .CK(n_120), .Q(\o_buffer[18] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][6]  (.D(n_132_310), .CK(n_120), .Q(\o_buffer[18] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][5]  (.D(n_132_309), .CK(n_120), .Q(\o_buffer[18] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][4]  (.D(n_132_308), .CK(n_120), .Q(\o_buffer[18] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][3]  (.D(n_132_307), .CK(n_120), .Q(\o_buffer[18] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][2]  (.D(n_132_306), .CK(n_120), .Q(\o_buffer[18] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][1]  (.D(n_132_305), .CK(n_120), .Q(\o_buffer[18] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[18][0]  (.D(n_132_304), .CK(n_120), .Q(\o_buffer[18] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][15]  (.D(n_132_303), .CK(n_120), .Q(
      \o_buffer[17] [15]), .QN());
   DFF_X1 \o_buffer_reg[17][14]  (.D(n_132_302), .CK(n_120), .Q(
      \o_buffer[17] [14]), .QN());
   DFF_X1 \o_buffer_reg[17][13]  (.D(n_132_301), .CK(n_120), .Q(
      \o_buffer[17] [13]), .QN());
   DFF_X1 \o_buffer_reg[17][12]  (.D(n_132_300), .CK(n_120), .Q(
      \o_buffer[17] [12]), .QN());
   DFF_X1 \o_buffer_reg[17][11]  (.D(n_132_299), .CK(n_120), .Q(
      \o_buffer[17] [11]), .QN());
   DFF_X1 \o_buffer_reg[17][10]  (.D(n_132_298), .CK(n_120), .Q(
      \o_buffer[17] [10]), .QN());
   DFF_X1 \o_buffer_reg[17][9]  (.D(n_132_297), .CK(n_120), .Q(\o_buffer[17] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][8]  (.D(n_132_296), .CK(n_120), .Q(\o_buffer[17] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][7]  (.D(n_132_295), .CK(n_120), .Q(\o_buffer[17] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][6]  (.D(n_132_294), .CK(n_120), .Q(\o_buffer[17] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][5]  (.D(n_132_293), .CK(n_120), .Q(\o_buffer[17] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][4]  (.D(n_132_292), .CK(n_120), .Q(\o_buffer[17] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][3]  (.D(n_132_291), .CK(n_120), .Q(\o_buffer[17] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][2]  (.D(n_132_290), .CK(n_120), .Q(\o_buffer[17] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][1]  (.D(n_132_289), .CK(n_120), .Q(\o_buffer[17] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[17][0]  (.D(n_132_288), .CK(n_120), .Q(\o_buffer[17] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][15]  (.D(n_132_287), .CK(n_120), .Q(
      \o_buffer[16] [15]), .QN());
   DFF_X1 \o_buffer_reg[16][14]  (.D(n_132_286), .CK(n_120), .Q(
      \o_buffer[16] [14]), .QN());
   DFF_X1 \o_buffer_reg[16][13]  (.D(n_132_285), .CK(n_120), .Q(
      \o_buffer[16] [13]), .QN());
   DFF_X1 \o_buffer_reg[16][12]  (.D(n_132_284), .CK(n_120), .Q(
      \o_buffer[16] [12]), .QN());
   DFF_X1 \o_buffer_reg[16][11]  (.D(n_132_283), .CK(n_120), .Q(
      \o_buffer[16] [11]), .QN());
   DFF_X1 \o_buffer_reg[16][10]  (.D(n_132_282), .CK(n_120), .Q(
      \o_buffer[16] [10]), .QN());
   DFF_X1 \o_buffer_reg[16][9]  (.D(n_132_281), .CK(n_120), .Q(\o_buffer[16] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][8]  (.D(n_132_280), .CK(n_120), .Q(\o_buffer[16] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][7]  (.D(n_132_279), .CK(n_120), .Q(\o_buffer[16] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][6]  (.D(n_132_278), .CK(n_120), .Q(\o_buffer[16] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][5]  (.D(n_132_277), .CK(n_120), .Q(\o_buffer[16] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][4]  (.D(n_132_276), .CK(n_120), .Q(\o_buffer[16] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][3]  (.D(n_132_275), .CK(n_120), .Q(\o_buffer[16] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][2]  (.D(n_132_274), .CK(n_120), .Q(\o_buffer[16] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][1]  (.D(n_132_273), .CK(n_120), .Q(\o_buffer[16] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[16][0]  (.D(n_132_272), .CK(n_120), .Q(\o_buffer[16] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][15]  (.D(n_132_271), .CK(n_120), .Q(
      \o_buffer[15] [15]), .QN());
   DFF_X1 \o_buffer_reg[15][14]  (.D(n_132_270), .CK(n_120), .Q(
      \o_buffer[15] [14]), .QN());
   DFF_X1 \o_buffer_reg[15][13]  (.D(n_132_269), .CK(n_120), .Q(
      \o_buffer[15] [13]), .QN());
   DFF_X1 \o_buffer_reg[15][12]  (.D(n_132_268), .CK(n_120), .Q(
      \o_buffer[15] [12]), .QN());
   DFF_X1 \o_buffer_reg[15][11]  (.D(n_132_267), .CK(n_120), .Q(
      \o_buffer[15] [11]), .QN());
   DFF_X1 \o_buffer_reg[15][10]  (.D(n_132_266), .CK(n_120), .Q(
      \o_buffer[15] [10]), .QN());
   DFF_X1 \o_buffer_reg[15][9]  (.D(n_132_265), .CK(n_120), .Q(\o_buffer[15] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][8]  (.D(n_132_264), .CK(n_120), .Q(\o_buffer[15] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][7]  (.D(n_132_263), .CK(n_120), .Q(\o_buffer[15] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][6]  (.D(n_132_262), .CK(n_120), .Q(\o_buffer[15] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][5]  (.D(n_132_261), .CK(n_120), .Q(\o_buffer[15] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][4]  (.D(n_132_260), .CK(n_120), .Q(\o_buffer[15] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][3]  (.D(n_132_259), .CK(n_120), .Q(\o_buffer[15] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][2]  (.D(n_132_258), .CK(n_120), .Q(\o_buffer[15] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][1]  (.D(n_132_257), .CK(n_120), .Q(\o_buffer[15] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[15][0]  (.D(n_132_256), .CK(n_120), .Q(\o_buffer[15] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][15]  (.D(n_132_255), .CK(n_120), .Q(
      \o_buffer[14] [15]), .QN());
   DFF_X1 \o_buffer_reg[14][14]  (.D(n_132_254), .CK(n_120), .Q(
      \o_buffer[14] [14]), .QN());
   DFF_X1 \o_buffer_reg[14][13]  (.D(n_132_253), .CK(n_120), .Q(
      \o_buffer[14] [13]), .QN());
   DFF_X1 \o_buffer_reg[14][12]  (.D(n_132_252), .CK(n_120), .Q(
      \o_buffer[14] [12]), .QN());
   DFF_X1 \o_buffer_reg[14][11]  (.D(n_132_251), .CK(n_120), .Q(
      \o_buffer[14] [11]), .QN());
   DFF_X1 \o_buffer_reg[14][10]  (.D(n_132_250), .CK(n_120), .Q(
      \o_buffer[14] [10]), .QN());
   DFF_X1 \o_buffer_reg[14][9]  (.D(n_132_249), .CK(n_120), .Q(\o_buffer[14] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][8]  (.D(n_132_248), .CK(n_120), .Q(\o_buffer[14] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][7]  (.D(n_132_247), .CK(n_120), .Q(\o_buffer[14] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][6]  (.D(n_132_246), .CK(n_120), .Q(\o_buffer[14] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][5]  (.D(n_132_245), .CK(n_120), .Q(\o_buffer[14] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][4]  (.D(n_132_244), .CK(n_120), .Q(\o_buffer[14] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][3]  (.D(n_132_243), .CK(n_120), .Q(\o_buffer[14] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][2]  (.D(n_132_242), .CK(n_120), .Q(\o_buffer[14] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][1]  (.D(n_132_241), .CK(n_120), .Q(\o_buffer[14] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[14][0]  (.D(n_132_240), .CK(n_120), .Q(\o_buffer[14] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][15]  (.D(n_132_239), .CK(n_120), .Q(
      \o_buffer[13] [15]), .QN());
   DFF_X1 \o_buffer_reg[13][14]  (.D(n_132_238), .CK(n_120), .Q(
      \o_buffer[13] [14]), .QN());
   DFF_X1 \o_buffer_reg[13][13]  (.D(n_132_237), .CK(n_120), .Q(
      \o_buffer[13] [13]), .QN());
   DFF_X1 \o_buffer_reg[13][12]  (.D(n_132_236), .CK(n_120), .Q(
      \o_buffer[13] [12]), .QN());
   DFF_X1 \o_buffer_reg[13][11]  (.D(n_132_235), .CK(n_120), .Q(
      \o_buffer[13] [11]), .QN());
   DFF_X1 \o_buffer_reg[13][10]  (.D(n_132_234), .CK(n_120), .Q(
      \o_buffer[13] [10]), .QN());
   DFF_X1 \o_buffer_reg[13][9]  (.D(n_132_233), .CK(n_120), .Q(\o_buffer[13] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][8]  (.D(n_132_232), .CK(n_120), .Q(\o_buffer[13] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][7]  (.D(n_132_231), .CK(n_120), .Q(\o_buffer[13] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][6]  (.D(n_132_230), .CK(n_120), .Q(\o_buffer[13] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][5]  (.D(n_132_229), .CK(n_120), .Q(\o_buffer[13] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][4]  (.D(n_132_228), .CK(n_120), .Q(\o_buffer[13] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][3]  (.D(n_132_227), .CK(n_120), .Q(\o_buffer[13] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][2]  (.D(n_132_226), .CK(n_120), .Q(\o_buffer[13] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][1]  (.D(n_132_225), .CK(n_120), .Q(\o_buffer[13] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[13][0]  (.D(n_132_224), .CK(n_120), .Q(\o_buffer[13] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][15]  (.D(n_132_223), .CK(n_120), .Q(
      \o_buffer[12] [15]), .QN());
   DFF_X1 \o_buffer_reg[12][14]  (.D(n_132_222), .CK(n_120), .Q(
      \o_buffer[12] [14]), .QN());
   DFF_X1 \o_buffer_reg[12][13]  (.D(n_132_221), .CK(n_120), .Q(
      \o_buffer[12] [13]), .QN());
   DFF_X1 \o_buffer_reg[12][12]  (.D(n_132_220), .CK(n_120), .Q(
      \o_buffer[12] [12]), .QN());
   DFF_X1 \o_buffer_reg[12][11]  (.D(n_132_219), .CK(n_120), .Q(
      \o_buffer[12] [11]), .QN());
   DFF_X1 \o_buffer_reg[12][10]  (.D(n_132_218), .CK(n_120), .Q(
      \o_buffer[12] [10]), .QN());
   DFF_X1 \o_buffer_reg[12][9]  (.D(n_132_217), .CK(n_120), .Q(\o_buffer[12] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][8]  (.D(n_132_216), .CK(n_120), .Q(\o_buffer[12] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][7]  (.D(n_132_215), .CK(n_120), .Q(\o_buffer[12] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][6]  (.D(n_132_214), .CK(n_120), .Q(\o_buffer[12] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][5]  (.D(n_132_213), .CK(n_120), .Q(\o_buffer[12] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][4]  (.D(n_132_212), .CK(n_120), .Q(\o_buffer[12] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][3]  (.D(n_132_211), .CK(n_120), .Q(\o_buffer[12] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][2]  (.D(n_132_210), .CK(n_120), .Q(\o_buffer[12] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][1]  (.D(n_132_209), .CK(n_120), .Q(\o_buffer[12] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[12][0]  (.D(n_132_208), .CK(n_120), .Q(\o_buffer[12] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][15]  (.D(n_132_207), .CK(n_120), .Q(
      \o_buffer[11] [15]), .QN());
   DFF_X1 \o_buffer_reg[11][14]  (.D(n_132_206), .CK(n_120), .Q(
      \o_buffer[11] [14]), .QN());
   DFF_X1 \o_buffer_reg[11][13]  (.D(n_132_205), .CK(n_120), .Q(
      \o_buffer[11] [13]), .QN());
   DFF_X1 \o_buffer_reg[11][12]  (.D(n_132_204), .CK(n_120), .Q(
      \o_buffer[11] [12]), .QN());
   DFF_X1 \o_buffer_reg[11][11]  (.D(n_132_203), .CK(n_120), .Q(
      \o_buffer[11] [11]), .QN());
   DFF_X1 \o_buffer_reg[11][10]  (.D(n_132_202), .CK(n_120), .Q(
      \o_buffer[11] [10]), .QN());
   DFF_X1 \o_buffer_reg[11][9]  (.D(n_132_201), .CK(n_120), .Q(\o_buffer[11] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][8]  (.D(n_132_200), .CK(n_120), .Q(\o_buffer[11] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][7]  (.D(n_132_199), .CK(n_120), .Q(\o_buffer[11] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][6]  (.D(n_132_198), .CK(n_120), .Q(\o_buffer[11] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][5]  (.D(n_132_197), .CK(n_120), .Q(\o_buffer[11] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][4]  (.D(n_132_196), .CK(n_120), .Q(\o_buffer[11] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][3]  (.D(n_132_195), .CK(n_120), .Q(\o_buffer[11] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][2]  (.D(n_132_194), .CK(n_120), .Q(\o_buffer[11] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][1]  (.D(n_132_193), .CK(n_120), .Q(\o_buffer[11] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[11][0]  (.D(n_132_192), .CK(n_120), .Q(\o_buffer[11] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][15]  (.D(n_132_191), .CK(n_120), .Q(
      \o_buffer[10] [15]), .QN());
   DFF_X1 \o_buffer_reg[10][14]  (.D(n_132_190), .CK(n_120), .Q(
      \o_buffer[10] [14]), .QN());
   DFF_X1 \o_buffer_reg[10][13]  (.D(n_132_189), .CK(n_120), .Q(
      \o_buffer[10] [13]), .QN());
   DFF_X1 \o_buffer_reg[10][12]  (.D(n_132_188), .CK(n_120), .Q(
      \o_buffer[10] [12]), .QN());
   DFF_X1 \o_buffer_reg[10][11]  (.D(n_132_187), .CK(n_120), .Q(
      \o_buffer[10] [11]), .QN());
   DFF_X1 \o_buffer_reg[10][10]  (.D(n_132_186), .CK(n_120), .Q(
      \o_buffer[10] [10]), .QN());
   DFF_X1 \o_buffer_reg[10][9]  (.D(n_132_185), .CK(n_120), .Q(\o_buffer[10] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][8]  (.D(n_132_184), .CK(n_120), .Q(\o_buffer[10] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][7]  (.D(n_132_183), .CK(n_120), .Q(\o_buffer[10] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][6]  (.D(n_132_182), .CK(n_120), .Q(\o_buffer[10] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][5]  (.D(n_132_181), .CK(n_120), .Q(\o_buffer[10] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][4]  (.D(n_132_180), .CK(n_120), .Q(\o_buffer[10] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][3]  (.D(n_132_179), .CK(n_120), .Q(\o_buffer[10] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][2]  (.D(n_132_178), .CK(n_120), .Q(\o_buffer[10] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][1]  (.D(n_132_177), .CK(n_120), .Q(\o_buffer[10] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[10][0]  (.D(n_132_176), .CK(n_120), .Q(\o_buffer[10] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][15]  (.D(n_132_175), .CK(n_120), .Q(\o_buffer[9] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][14]  (.D(n_132_174), .CK(n_120), .Q(\o_buffer[9] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][13]  (.D(n_132_173), .CK(n_120), .Q(\o_buffer[9] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][12]  (.D(n_132_172), .CK(n_120), .Q(\o_buffer[9] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][11]  (.D(n_132_171), .CK(n_120), .Q(\o_buffer[9] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][10]  (.D(n_132_170), .CK(n_120), .Q(\o_buffer[9] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][9]  (.D(n_132_169), .CK(n_120), .Q(\o_buffer[9] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][8]  (.D(n_132_168), .CK(n_120), .Q(\o_buffer[9] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][7]  (.D(n_132_167), .CK(n_120), .Q(\o_buffer[9] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][6]  (.D(n_132_166), .CK(n_120), .Q(\o_buffer[9] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][5]  (.D(n_132_165), .CK(n_120), .Q(\o_buffer[9] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][4]  (.D(n_132_164), .CK(n_120), .Q(\o_buffer[9] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][3]  (.D(n_132_163), .CK(n_120), .Q(\o_buffer[9] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][2]  (.D(n_132_162), .CK(n_120), .Q(\o_buffer[9] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][1]  (.D(n_132_161), .CK(n_120), .Q(\o_buffer[9] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[9][0]  (.D(n_132_160), .CK(n_120), .Q(\o_buffer[9] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][15]  (.D(n_132_159), .CK(n_120), .Q(\o_buffer[8] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][14]  (.D(n_132_158), .CK(n_120), .Q(\o_buffer[8] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][13]  (.D(n_132_157), .CK(n_120), .Q(\o_buffer[8] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][12]  (.D(n_132_156), .CK(n_120), .Q(\o_buffer[8] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][11]  (.D(n_132_155), .CK(n_120), .Q(\o_buffer[8] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][10]  (.D(n_132_154), .CK(n_120), .Q(\o_buffer[8] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][9]  (.D(n_132_153), .CK(n_120), .Q(\o_buffer[8] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][8]  (.D(n_132_152), .CK(n_120), .Q(\o_buffer[8] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][7]  (.D(n_132_151), .CK(n_120), .Q(\o_buffer[8] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][6]  (.D(n_132_150), .CK(n_120), .Q(\o_buffer[8] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][5]  (.D(n_132_149), .CK(n_120), .Q(\o_buffer[8] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][4]  (.D(n_132_148), .CK(n_120), .Q(\o_buffer[8] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][3]  (.D(n_132_147), .CK(n_120), .Q(\o_buffer[8] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][2]  (.D(n_132_146), .CK(n_120), .Q(\o_buffer[8] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][1]  (.D(n_132_145), .CK(n_120), .Q(\o_buffer[8] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[8][0]  (.D(n_132_144), .CK(n_120), .Q(\o_buffer[8] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][15]  (.D(n_132_143), .CK(n_120), .Q(\o_buffer[7] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][14]  (.D(n_132_142), .CK(n_120), .Q(\o_buffer[7] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][13]  (.D(n_132_141), .CK(n_120), .Q(\o_buffer[7] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][12]  (.D(n_132_140), .CK(n_120), .Q(\o_buffer[7] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][11]  (.D(n_132_139), .CK(n_120), .Q(\o_buffer[7] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][10]  (.D(n_132_138), .CK(n_120), .Q(\o_buffer[7] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][9]  (.D(n_132_137), .CK(n_120), .Q(\o_buffer[7] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][8]  (.D(n_132_136), .CK(n_120), .Q(\o_buffer[7] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][7]  (.D(n_132_135), .CK(n_120), .Q(\o_buffer[7] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][6]  (.D(n_132_134), .CK(n_120), .Q(\o_buffer[7] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][5]  (.D(n_132_133), .CK(n_120), .Q(\o_buffer[7] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][4]  (.D(n_132_132), .CK(n_120), .Q(\o_buffer[7] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][3]  (.D(n_132_131), .CK(n_120), .Q(\o_buffer[7] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][2]  (.D(n_132_130), .CK(n_120), .Q(\o_buffer[7] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][1]  (.D(n_132_129), .CK(n_120), .Q(\o_buffer[7] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[7][0]  (.D(n_132_128), .CK(n_120), .Q(\o_buffer[7] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][15]  (.D(n_132_127), .CK(n_120), .Q(\o_buffer[6] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][14]  (.D(n_132_126), .CK(n_120), .Q(\o_buffer[6] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][13]  (.D(n_132_125), .CK(n_120), .Q(\o_buffer[6] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][12]  (.D(n_132_124), .CK(n_120), .Q(\o_buffer[6] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][11]  (.D(n_132_123), .CK(n_120), .Q(\o_buffer[6] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][10]  (.D(n_132_122), .CK(n_120), .Q(\o_buffer[6] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][9]  (.D(n_132_121), .CK(n_120), .Q(\o_buffer[6] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][8]  (.D(n_132_120), .CK(n_120), .Q(\o_buffer[6] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][7]  (.D(n_132_119), .CK(n_120), .Q(\o_buffer[6] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][6]  (.D(n_132_118), .CK(n_120), .Q(\o_buffer[6] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][5]  (.D(n_132_117), .CK(n_120), .Q(\o_buffer[6] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][4]  (.D(n_132_116), .CK(n_120), .Q(\o_buffer[6] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][3]  (.D(n_132_115), .CK(n_120), .Q(\o_buffer[6] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][2]  (.D(n_132_114), .CK(n_120), .Q(\o_buffer[6] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][1]  (.D(n_132_113), .CK(n_120), .Q(\o_buffer[6] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[6][0]  (.D(n_132_112), .CK(n_120), .Q(\o_buffer[6] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][15]  (.D(n_132_111), .CK(n_120), .Q(\o_buffer[5] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][14]  (.D(n_132_110), .CK(n_120), .Q(\o_buffer[5] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][13]  (.D(n_132_109), .CK(n_120), .Q(\o_buffer[5] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][12]  (.D(n_132_108), .CK(n_120), .Q(\o_buffer[5] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][11]  (.D(n_132_107), .CK(n_120), .Q(\o_buffer[5] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][10]  (.D(n_132_106), .CK(n_120), .Q(\o_buffer[5] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][9]  (.D(n_132_105), .CK(n_120), .Q(\o_buffer[5] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][8]  (.D(n_132_104), .CK(n_120), .Q(\o_buffer[5] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][7]  (.D(n_132_103), .CK(n_120), .Q(\o_buffer[5] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][6]  (.D(n_132_102), .CK(n_120), .Q(\o_buffer[5] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][5]  (.D(n_132_101), .CK(n_120), .Q(\o_buffer[5] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][4]  (.D(n_132_100), .CK(n_120), .Q(\o_buffer[5] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][3]  (.D(n_132_99), .CK(n_120), .Q(\o_buffer[5] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][2]  (.D(n_132_98), .CK(n_120), .Q(\o_buffer[5] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][1]  (.D(n_132_97), .CK(n_120), .Q(\o_buffer[5] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[5][0]  (.D(n_132_96), .CK(n_120), .Q(\o_buffer[5] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][15]  (.D(n_132_95), .CK(n_120), .Q(\o_buffer[4] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][14]  (.D(n_132_94), .CK(n_120), .Q(\o_buffer[4] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][13]  (.D(n_132_93), .CK(n_120), .Q(\o_buffer[4] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][12]  (.D(n_132_92), .CK(n_120), .Q(\o_buffer[4] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][11]  (.D(n_132_91), .CK(n_120), .Q(\o_buffer[4] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][10]  (.D(n_132_90), .CK(n_120), .Q(\o_buffer[4] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][9]  (.D(n_132_89), .CK(n_120), .Q(\o_buffer[4] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][8]  (.D(n_132_88), .CK(n_120), .Q(\o_buffer[4] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][7]  (.D(n_132_87), .CK(n_120), .Q(\o_buffer[4] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][6]  (.D(n_132_86), .CK(n_120), .Q(\o_buffer[4] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][5]  (.D(n_132_85), .CK(n_120), .Q(\o_buffer[4] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][4]  (.D(n_132_84), .CK(n_120), .Q(\o_buffer[4] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][3]  (.D(n_132_83), .CK(n_120), .Q(\o_buffer[4] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][2]  (.D(n_132_82), .CK(n_120), .Q(\o_buffer[4] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][1]  (.D(n_132_81), .CK(n_120), .Q(\o_buffer[4] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[4][0]  (.D(n_132_80), .CK(n_120), .Q(\o_buffer[4] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][15]  (.D(n_132_79), .CK(n_120), .Q(\o_buffer[3] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][14]  (.D(n_132_78), .CK(n_120), .Q(\o_buffer[3] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][13]  (.D(n_132_77), .CK(n_120), .Q(\o_buffer[3] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][12]  (.D(n_132_76), .CK(n_120), .Q(\o_buffer[3] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][11]  (.D(n_132_75), .CK(n_120), .Q(\o_buffer[3] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][10]  (.D(n_132_74), .CK(n_120), .Q(\o_buffer[3] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][9]  (.D(n_132_73), .CK(n_120), .Q(\o_buffer[3] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][8]  (.D(n_132_72), .CK(n_120), .Q(\o_buffer[3] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][7]  (.D(n_132_71), .CK(n_120), .Q(\o_buffer[3] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][6]  (.D(n_132_70), .CK(n_120), .Q(\o_buffer[3] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][5]  (.D(n_132_69), .CK(n_120), .Q(\o_buffer[3] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][4]  (.D(n_132_68), .CK(n_120), .Q(\o_buffer[3] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][3]  (.D(n_132_67), .CK(n_120), .Q(\o_buffer[3] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][2]  (.D(n_132_66), .CK(n_120), .Q(\o_buffer[3] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][1]  (.D(n_132_65), .CK(n_120), .Q(\o_buffer[3] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[3][0]  (.D(n_132_64), .CK(n_120), .Q(\o_buffer[3] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][15]  (.D(n_132_63), .CK(n_120), .Q(\o_buffer[2] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][14]  (.D(n_132_62), .CK(n_120), .Q(\o_buffer[2] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][13]  (.D(n_132_61), .CK(n_120), .Q(\o_buffer[2] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][12]  (.D(n_132_60), .CK(n_120), .Q(\o_buffer[2] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][11]  (.D(n_132_59), .CK(n_120), .Q(\o_buffer[2] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][10]  (.D(n_132_58), .CK(n_120), .Q(\o_buffer[2] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][9]  (.D(n_132_57), .CK(n_120), .Q(\o_buffer[2] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][8]  (.D(n_132_56), .CK(n_120), .Q(\o_buffer[2] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][7]  (.D(n_132_55), .CK(n_120), .Q(\o_buffer[2] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][6]  (.D(n_132_54), .CK(n_120), .Q(\o_buffer[2] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][5]  (.D(n_132_53), .CK(n_120), .Q(\o_buffer[2] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][4]  (.D(n_132_52), .CK(n_120), .Q(\o_buffer[2] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][3]  (.D(n_132_51), .CK(n_120), .Q(\o_buffer[2] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][2]  (.D(n_132_50), .CK(n_120), .Q(\o_buffer[2] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][1]  (.D(n_132_49), .CK(n_120), .Q(\o_buffer[2] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[2][0]  (.D(n_132_48), .CK(n_120), .Q(\o_buffer[2] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][15]  (.D(n_132_47), .CK(n_120), .Q(\o_buffer[1] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][14]  (.D(n_132_46), .CK(n_120), .Q(\o_buffer[1] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][13]  (.D(n_132_45), .CK(n_120), .Q(\o_buffer[1] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][12]  (.D(n_132_44), .CK(n_120), .Q(\o_buffer[1] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][11]  (.D(n_132_43), .CK(n_120), .Q(\o_buffer[1] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][10]  (.D(n_132_42), .CK(n_120), .Q(\o_buffer[1] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][9]  (.D(n_132_41), .CK(n_120), .Q(\o_buffer[1] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][8]  (.D(n_132_40), .CK(n_120), .Q(\o_buffer[1] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][7]  (.D(n_132_39), .CK(n_120), .Q(\o_buffer[1] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][6]  (.D(n_132_38), .CK(n_120), .Q(\o_buffer[1] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][5]  (.D(n_132_37), .CK(n_120), .Q(\o_buffer[1] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][4]  (.D(n_132_36), .CK(n_120), .Q(\o_buffer[1] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][3]  (.D(n_132_35), .CK(n_120), .Q(\o_buffer[1] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][2]  (.D(n_132_34), .CK(n_120), .Q(\o_buffer[1] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][1]  (.D(n_132_33), .CK(n_120), .Q(\o_buffer[1] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[1][0]  (.D(n_132_32), .CK(n_120), .Q(\o_buffer[1] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][15]  (.D(n_132_31), .CK(n_120), .Q(\o_buffer[0] [15]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][14]  (.D(n_132_30), .CK(n_120), .Q(\o_buffer[0] [14]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][13]  (.D(n_132_29), .CK(n_120), .Q(\o_buffer[0] [13]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][12]  (.D(n_132_28), .CK(n_120), .Q(\o_buffer[0] [12]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][11]  (.D(n_132_27), .CK(n_120), .Q(\o_buffer[0] [11]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][10]  (.D(n_132_26), .CK(n_120), .Q(\o_buffer[0] [10]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][9]  (.D(n_132_25), .CK(n_120), .Q(\o_buffer[0] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][8]  (.D(n_132_24), .CK(n_120), .Q(\o_buffer[0] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][7]  (.D(n_132_23), .CK(n_120), .Q(\o_buffer[0] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][6]  (.D(n_132_22), .CK(n_120), .Q(\o_buffer[0] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][5]  (.D(n_132_21), .CK(n_120), .Q(\o_buffer[0] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][4]  (.D(n_132_20), .CK(n_120), .Q(\o_buffer[0] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][3]  (.D(n_132_19), .CK(n_120), .Q(\o_buffer[0] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][2]  (.D(n_132_18), .CK(n_120), .Q(\o_buffer[0] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][1]  (.D(n_132_17), .CK(n_120), .Q(\o_buffer[0] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[0][0]  (.D(n_132_16), .CK(n_120), .Q(\o_buffer[0] [0]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][15]  (.D(n_132_15), .CK(n_120), .Q(
      \o_buffer[119] [15]), .QN());
   DFF_X1 \o_buffer_reg[119][14]  (.D(n_132_14), .CK(n_120), .Q(
      \o_buffer[119] [14]), .QN());
   DFF_X1 \o_buffer_reg[119][13]  (.D(n_132_13), .CK(n_120), .Q(
      \o_buffer[119] [13]), .QN());
   DFF_X1 \o_buffer_reg[119][12]  (.D(n_132_12), .CK(n_120), .Q(
      \o_buffer[119] [12]), .QN());
   DFF_X1 \o_buffer_reg[119][11]  (.D(n_132_11), .CK(n_120), .Q(
      \o_buffer[119] [11]), .QN());
   DFF_X1 \o_buffer_reg[119][10]  (.D(n_132_10), .CK(n_120), .Q(
      \o_buffer[119] [10]), .QN());
   DFF_X1 \o_buffer_reg[119][9]  (.D(n_132_9), .CK(n_120), .Q(\o_buffer[119] [9]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][8]  (.D(n_132_8), .CK(n_120), .Q(\o_buffer[119] [8]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][7]  (.D(n_132_7), .CK(n_120), .Q(\o_buffer[119] [7]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][6]  (.D(n_132_6), .CK(n_120), .Q(\o_buffer[119] [6]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][5]  (.D(n_132_5), .CK(n_120), .Q(\o_buffer[119] [5]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][4]  (.D(n_132_4), .CK(n_120), .Q(\o_buffer[119] [4]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][3]  (.D(n_132_3), .CK(n_120), .Q(\o_buffer[119] [3]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][2]  (.D(n_132_2), .CK(n_120), .Q(\o_buffer[119] [2]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][1]  (.D(n_132_1), .CK(n_120), .Q(\o_buffer[119] [1]), 
      .QN());
   DFF_X1 \o_buffer_reg[119][0]  (.D(n_132_0), .CK(n_120), .Q(\o_buffer[119] [0]), 
      .QN());
   MUX2_X1 i_132_0_0 (.A(\o_buffer[58] [15]), .B(i_mem_data[15]), .S(n_61), 
      .Z(n_132_959));
   MUX2_X1 i_132_0_1 (.A(\o_buffer[58] [14]), .B(i_mem_data[14]), .S(n_61), 
      .Z(n_132_958));
   MUX2_X1 i_132_0_2 (.A(\o_buffer[58] [13]), .B(i_mem_data[13]), .S(n_61), 
      .Z(n_132_957));
   MUX2_X1 i_132_0_3 (.A(\o_buffer[58] [12]), .B(i_mem_data[12]), .S(n_61), 
      .Z(n_132_956));
   MUX2_X1 i_132_0_4 (.A(\o_buffer[58] [11]), .B(i_mem_data[11]), .S(n_61), 
      .Z(n_132_955));
   MUX2_X1 i_132_0_5 (.A(\o_buffer[58] [10]), .B(i_mem_data[10]), .S(n_61), 
      .Z(n_132_954));
   MUX2_X1 i_132_0_6 (.A(\o_buffer[58] [9]), .B(i_mem_data[9]), .S(n_61), 
      .Z(n_132_953));
   MUX2_X1 i_132_0_7 (.A(\o_buffer[58] [8]), .B(i_mem_data[8]), .S(n_61), 
      .Z(n_132_952));
   MUX2_X1 i_132_0_8 (.A(\o_buffer[58] [7]), .B(i_mem_data[7]), .S(n_61), 
      .Z(n_132_951));
   MUX2_X1 i_132_0_9 (.A(\o_buffer[58] [6]), .B(i_mem_data[6]), .S(n_61), 
      .Z(n_132_950));
   MUX2_X1 i_132_0_10 (.A(\o_buffer[58] [5]), .B(i_mem_data[5]), .S(n_61), 
      .Z(n_132_949));
   MUX2_X1 i_132_0_11 (.A(\o_buffer[58] [4]), .B(i_mem_data[4]), .S(n_61), 
      .Z(n_132_948));
   MUX2_X1 i_132_0_12 (.A(\o_buffer[58] [3]), .B(i_mem_data[3]), .S(n_61), 
      .Z(n_132_947));
   MUX2_X1 i_132_0_13 (.A(\o_buffer[58] [2]), .B(i_mem_data[2]), .S(n_61), 
      .Z(n_132_946));
   MUX2_X1 i_132_0_14 (.A(\o_buffer[58] [1]), .B(i_mem_data[1]), .S(n_61), 
      .Z(n_132_945));
   MUX2_X1 i_132_0_15 (.A(\o_buffer[58] [0]), .B(i_mem_data[0]), .S(n_61), 
      .Z(n_132_944));
   MUX2_X1 i_132_0_16 (.A(\o_buffer[57] [15]), .B(i_mem_data[15]), .S(n_62), 
      .Z(n_132_943));
   MUX2_X1 i_132_0_17 (.A(\o_buffer[57] [14]), .B(i_mem_data[14]), .S(n_62), 
      .Z(n_132_942));
   MUX2_X1 i_132_0_18 (.A(\o_buffer[57] [13]), .B(i_mem_data[13]), .S(n_62), 
      .Z(n_132_941));
   MUX2_X1 i_132_0_19 (.A(\o_buffer[57] [12]), .B(i_mem_data[12]), .S(n_62), 
      .Z(n_132_940));
   MUX2_X1 i_132_0_20 (.A(\o_buffer[57] [11]), .B(i_mem_data[11]), .S(n_62), 
      .Z(n_132_939));
   MUX2_X1 i_132_0_21 (.A(\o_buffer[57] [10]), .B(i_mem_data[10]), .S(n_62), 
      .Z(n_132_938));
   MUX2_X1 i_132_0_22 (.A(\o_buffer[57] [9]), .B(i_mem_data[9]), .S(n_62), 
      .Z(n_132_937));
   MUX2_X1 i_132_0_23 (.A(\o_buffer[57] [8]), .B(i_mem_data[8]), .S(n_62), 
      .Z(n_132_936));
   MUX2_X1 i_132_0_24 (.A(\o_buffer[57] [7]), .B(i_mem_data[7]), .S(n_62), 
      .Z(n_132_935));
   MUX2_X1 i_132_0_25 (.A(\o_buffer[57] [6]), .B(i_mem_data[6]), .S(n_62), 
      .Z(n_132_934));
   MUX2_X1 i_132_0_26 (.A(\o_buffer[57] [5]), .B(i_mem_data[5]), .S(n_62), 
      .Z(n_132_933));
   MUX2_X1 i_132_0_27 (.A(\o_buffer[57] [4]), .B(i_mem_data[4]), .S(n_62), 
      .Z(n_132_932));
   MUX2_X1 i_132_0_28 (.A(\o_buffer[57] [3]), .B(i_mem_data[3]), .S(n_62), 
      .Z(n_132_931));
   MUX2_X1 i_132_0_29 (.A(\o_buffer[57] [2]), .B(i_mem_data[2]), .S(n_62), 
      .Z(n_132_930));
   MUX2_X1 i_132_0_30 (.A(\o_buffer[57] [1]), .B(i_mem_data[1]), .S(n_62), 
      .Z(n_132_929));
   MUX2_X1 i_132_0_31 (.A(\o_buffer[57] [0]), .B(i_mem_data[0]), .S(n_62), 
      .Z(n_132_928));
   MUX2_X1 i_132_0_32 (.A(\o_buffer[56] [15]), .B(i_mem_data[15]), .S(n_63), 
      .Z(n_132_927));
   MUX2_X1 i_132_0_33 (.A(\o_buffer[56] [14]), .B(i_mem_data[14]), .S(n_63), 
      .Z(n_132_926));
   MUX2_X1 i_132_0_34 (.A(\o_buffer[56] [13]), .B(i_mem_data[13]), .S(n_63), 
      .Z(n_132_925));
   MUX2_X1 i_132_0_35 (.A(\o_buffer[56] [12]), .B(i_mem_data[12]), .S(n_63), 
      .Z(n_132_924));
   MUX2_X1 i_132_0_36 (.A(\o_buffer[56] [11]), .B(i_mem_data[11]), .S(n_63), 
      .Z(n_132_923));
   MUX2_X1 i_132_0_37 (.A(\o_buffer[56] [10]), .B(i_mem_data[10]), .S(n_63), 
      .Z(n_132_922));
   MUX2_X1 i_132_0_38 (.A(\o_buffer[56] [9]), .B(i_mem_data[9]), .S(n_63), 
      .Z(n_132_921));
   MUX2_X1 i_132_0_39 (.A(\o_buffer[56] [8]), .B(i_mem_data[8]), .S(n_63), 
      .Z(n_132_920));
   MUX2_X1 i_132_0_40 (.A(\o_buffer[56] [7]), .B(i_mem_data[7]), .S(n_63), 
      .Z(n_132_919));
   MUX2_X1 i_132_0_41 (.A(\o_buffer[56] [6]), .B(i_mem_data[6]), .S(n_63), 
      .Z(n_132_918));
   MUX2_X1 i_132_0_42 (.A(\o_buffer[56] [5]), .B(i_mem_data[5]), .S(n_63), 
      .Z(n_132_917));
   MUX2_X1 i_132_0_43 (.A(\o_buffer[56] [4]), .B(i_mem_data[4]), .S(n_63), 
      .Z(n_132_916));
   MUX2_X1 i_132_0_44 (.A(\o_buffer[56] [3]), .B(i_mem_data[3]), .S(n_63), 
      .Z(n_132_915));
   MUX2_X1 i_132_0_45 (.A(\o_buffer[56] [2]), .B(i_mem_data[2]), .S(n_63), 
      .Z(n_132_914));
   MUX2_X1 i_132_0_46 (.A(\o_buffer[56] [1]), .B(i_mem_data[1]), .S(n_63), 
      .Z(n_132_913));
   MUX2_X1 i_132_0_47 (.A(\o_buffer[56] [0]), .B(i_mem_data[0]), .S(n_63), 
      .Z(n_132_912));
   MUX2_X1 i_132_0_48 (.A(\o_buffer[55] [15]), .B(i_mem_data[15]), .S(n_64), 
      .Z(n_132_911));
   MUX2_X1 i_132_0_49 (.A(\o_buffer[55] [14]), .B(i_mem_data[14]), .S(n_64), 
      .Z(n_132_910));
   MUX2_X1 i_132_0_50 (.A(\o_buffer[55] [13]), .B(i_mem_data[13]), .S(n_64), 
      .Z(n_132_909));
   MUX2_X1 i_132_0_51 (.A(\o_buffer[55] [12]), .B(i_mem_data[12]), .S(n_64), 
      .Z(n_132_908));
   MUX2_X1 i_132_0_52 (.A(\o_buffer[55] [11]), .B(i_mem_data[11]), .S(n_64), 
      .Z(n_132_907));
   MUX2_X1 i_132_0_53 (.A(\o_buffer[55] [10]), .B(i_mem_data[10]), .S(n_64), 
      .Z(n_132_906));
   MUX2_X1 i_132_0_54 (.A(\o_buffer[55] [9]), .B(i_mem_data[9]), .S(n_64), 
      .Z(n_132_905));
   MUX2_X1 i_132_0_55 (.A(\o_buffer[55] [8]), .B(i_mem_data[8]), .S(n_64), 
      .Z(n_132_904));
   MUX2_X1 i_132_0_56 (.A(\o_buffer[55] [7]), .B(i_mem_data[7]), .S(n_64), 
      .Z(n_132_903));
   MUX2_X1 i_132_0_57 (.A(\o_buffer[55] [6]), .B(i_mem_data[6]), .S(n_64), 
      .Z(n_132_902));
   MUX2_X1 i_132_0_58 (.A(\o_buffer[55] [5]), .B(i_mem_data[5]), .S(n_64), 
      .Z(n_132_901));
   MUX2_X1 i_132_0_59 (.A(\o_buffer[55] [4]), .B(i_mem_data[4]), .S(n_64), 
      .Z(n_132_900));
   MUX2_X1 i_132_0_60 (.A(\o_buffer[55] [3]), .B(i_mem_data[3]), .S(n_64), 
      .Z(n_132_899));
   MUX2_X1 i_132_0_61 (.A(\o_buffer[55] [2]), .B(i_mem_data[2]), .S(n_64), 
      .Z(n_132_898));
   MUX2_X1 i_132_0_62 (.A(\o_buffer[55] [1]), .B(i_mem_data[1]), .S(n_64), 
      .Z(n_132_897));
   MUX2_X1 i_132_0_63 (.A(\o_buffer[55] [0]), .B(i_mem_data[0]), .S(n_64), 
      .Z(n_132_896));
   MUX2_X1 i_132_0_64 (.A(\o_buffer[54] [15]), .B(i_mem_data[15]), .S(n_65), 
      .Z(n_132_895));
   MUX2_X1 i_132_0_65 (.A(\o_buffer[54] [14]), .B(i_mem_data[14]), .S(n_65), 
      .Z(n_132_894));
   MUX2_X1 i_132_0_66 (.A(\o_buffer[54] [13]), .B(i_mem_data[13]), .S(n_65), 
      .Z(n_132_893));
   MUX2_X1 i_132_0_67 (.A(\o_buffer[54] [12]), .B(i_mem_data[12]), .S(n_65), 
      .Z(n_132_892));
   MUX2_X1 i_132_0_68 (.A(\o_buffer[54] [11]), .B(i_mem_data[11]), .S(n_65), 
      .Z(n_132_891));
   MUX2_X1 i_132_0_69 (.A(\o_buffer[54] [10]), .B(i_mem_data[10]), .S(n_65), 
      .Z(n_132_890));
   MUX2_X1 i_132_0_70 (.A(\o_buffer[54] [9]), .B(i_mem_data[9]), .S(n_65), 
      .Z(n_132_889));
   MUX2_X1 i_132_0_71 (.A(\o_buffer[54] [8]), .B(i_mem_data[8]), .S(n_65), 
      .Z(n_132_888));
   MUX2_X1 i_132_0_72 (.A(\o_buffer[54] [7]), .B(i_mem_data[7]), .S(n_65), 
      .Z(n_132_887));
   MUX2_X1 i_132_0_73 (.A(\o_buffer[54] [6]), .B(i_mem_data[6]), .S(n_65), 
      .Z(n_132_886));
   MUX2_X1 i_132_0_74 (.A(\o_buffer[54] [5]), .B(i_mem_data[5]), .S(n_65), 
      .Z(n_132_885));
   MUX2_X1 i_132_0_75 (.A(\o_buffer[54] [4]), .B(i_mem_data[4]), .S(n_65), 
      .Z(n_132_884));
   MUX2_X1 i_132_0_76 (.A(\o_buffer[54] [3]), .B(i_mem_data[3]), .S(n_65), 
      .Z(n_132_883));
   MUX2_X1 i_132_0_77 (.A(\o_buffer[54] [2]), .B(i_mem_data[2]), .S(n_65), 
      .Z(n_132_882));
   MUX2_X1 i_132_0_78 (.A(\o_buffer[54] [1]), .B(i_mem_data[1]), .S(n_65), 
      .Z(n_132_881));
   MUX2_X1 i_132_0_79 (.A(\o_buffer[54] [0]), .B(i_mem_data[0]), .S(n_65), 
      .Z(n_132_880));
   MUX2_X1 i_132_0_80 (.A(\o_buffer[53] [15]), .B(i_mem_data[15]), .S(n_66), 
      .Z(n_132_879));
   MUX2_X1 i_132_0_81 (.A(\o_buffer[53] [14]), .B(i_mem_data[14]), .S(n_66), 
      .Z(n_132_878));
   MUX2_X1 i_132_0_82 (.A(\o_buffer[53] [13]), .B(i_mem_data[13]), .S(n_66), 
      .Z(n_132_877));
   MUX2_X1 i_132_0_83 (.A(\o_buffer[53] [12]), .B(i_mem_data[12]), .S(n_66), 
      .Z(n_132_876));
   MUX2_X1 i_132_0_84 (.A(\o_buffer[53] [11]), .B(i_mem_data[11]), .S(n_66), 
      .Z(n_132_875));
   MUX2_X1 i_132_0_85 (.A(\o_buffer[53] [10]), .B(i_mem_data[10]), .S(n_66), 
      .Z(n_132_874));
   MUX2_X1 i_132_0_86 (.A(\o_buffer[53] [9]), .B(i_mem_data[9]), .S(n_66), 
      .Z(n_132_873));
   MUX2_X1 i_132_0_87 (.A(\o_buffer[53] [8]), .B(i_mem_data[8]), .S(n_66), 
      .Z(n_132_872));
   MUX2_X1 i_132_0_88 (.A(\o_buffer[53] [7]), .B(i_mem_data[7]), .S(n_66), 
      .Z(n_132_871));
   MUX2_X1 i_132_0_89 (.A(\o_buffer[53] [6]), .B(i_mem_data[6]), .S(n_66), 
      .Z(n_132_870));
   MUX2_X1 i_132_0_90 (.A(\o_buffer[53] [5]), .B(i_mem_data[5]), .S(n_66), 
      .Z(n_132_869));
   MUX2_X1 i_132_0_91 (.A(\o_buffer[53] [4]), .B(i_mem_data[4]), .S(n_66), 
      .Z(n_132_868));
   MUX2_X1 i_132_0_92 (.A(\o_buffer[53] [3]), .B(i_mem_data[3]), .S(n_66), 
      .Z(n_132_867));
   MUX2_X1 i_132_0_93 (.A(\o_buffer[53] [2]), .B(i_mem_data[2]), .S(n_66), 
      .Z(n_132_866));
   MUX2_X1 i_132_0_94 (.A(\o_buffer[53] [1]), .B(i_mem_data[1]), .S(n_66), 
      .Z(n_132_865));
   MUX2_X1 i_132_0_95 (.A(\o_buffer[53] [0]), .B(i_mem_data[0]), .S(n_66), 
      .Z(n_132_864));
   MUX2_X1 i_132_0_96 (.A(\o_buffer[52] [15]), .B(i_mem_data[15]), .S(n_67), 
      .Z(n_132_863));
   MUX2_X1 i_132_0_97 (.A(\o_buffer[52] [14]), .B(i_mem_data[14]), .S(n_67), 
      .Z(n_132_862));
   MUX2_X1 i_132_0_98 (.A(\o_buffer[52] [13]), .B(i_mem_data[13]), .S(n_67), 
      .Z(n_132_861));
   MUX2_X1 i_132_0_99 (.A(\o_buffer[52] [12]), .B(i_mem_data[12]), .S(n_67), 
      .Z(n_132_860));
   MUX2_X1 i_132_0_100 (.A(\o_buffer[52] [11]), .B(i_mem_data[11]), .S(n_67), 
      .Z(n_132_859));
   MUX2_X1 i_132_0_101 (.A(\o_buffer[52] [10]), .B(i_mem_data[10]), .S(n_67), 
      .Z(n_132_858));
   MUX2_X1 i_132_0_102 (.A(\o_buffer[52] [9]), .B(i_mem_data[9]), .S(n_67), 
      .Z(n_132_857));
   MUX2_X1 i_132_0_103 (.A(\o_buffer[52] [8]), .B(i_mem_data[8]), .S(n_67), 
      .Z(n_132_856));
   MUX2_X1 i_132_0_104 (.A(\o_buffer[52] [7]), .B(i_mem_data[7]), .S(n_67), 
      .Z(n_132_855));
   MUX2_X1 i_132_0_105 (.A(\o_buffer[52] [6]), .B(i_mem_data[6]), .S(n_67), 
      .Z(n_132_854));
   MUX2_X1 i_132_0_106 (.A(\o_buffer[52] [5]), .B(i_mem_data[5]), .S(n_67), 
      .Z(n_132_853));
   MUX2_X1 i_132_0_107 (.A(\o_buffer[52] [4]), .B(i_mem_data[4]), .S(n_67), 
      .Z(n_132_852));
   MUX2_X1 i_132_0_108 (.A(\o_buffer[52] [3]), .B(i_mem_data[3]), .S(n_67), 
      .Z(n_132_851));
   MUX2_X1 i_132_0_109 (.A(\o_buffer[52] [2]), .B(i_mem_data[2]), .S(n_67), 
      .Z(n_132_850));
   MUX2_X1 i_132_0_110 (.A(\o_buffer[52] [1]), .B(i_mem_data[1]), .S(n_67), 
      .Z(n_132_849));
   MUX2_X1 i_132_0_111 (.A(\o_buffer[52] [0]), .B(i_mem_data[0]), .S(n_67), 
      .Z(n_132_848));
   MUX2_X1 i_132_0_112 (.A(\o_buffer[51] [15]), .B(i_mem_data[15]), .S(n_68), 
      .Z(n_132_847));
   MUX2_X1 i_132_0_113 (.A(\o_buffer[51] [14]), .B(i_mem_data[14]), .S(n_68), 
      .Z(n_132_846));
   MUX2_X1 i_132_0_114 (.A(\o_buffer[51] [13]), .B(i_mem_data[13]), .S(n_68), 
      .Z(n_132_845));
   MUX2_X1 i_132_0_115 (.A(\o_buffer[51] [12]), .B(i_mem_data[12]), .S(n_68), 
      .Z(n_132_844));
   MUX2_X1 i_132_0_116 (.A(\o_buffer[51] [11]), .B(i_mem_data[11]), .S(n_68), 
      .Z(n_132_843));
   MUX2_X1 i_132_0_117 (.A(\o_buffer[51] [10]), .B(i_mem_data[10]), .S(n_68), 
      .Z(n_132_842));
   MUX2_X1 i_132_0_118 (.A(\o_buffer[51] [9]), .B(i_mem_data[9]), .S(n_68), 
      .Z(n_132_841));
   MUX2_X1 i_132_0_119 (.A(\o_buffer[51] [8]), .B(i_mem_data[8]), .S(n_68), 
      .Z(n_132_840));
   MUX2_X1 i_132_0_120 (.A(\o_buffer[51] [7]), .B(i_mem_data[7]), .S(n_68), 
      .Z(n_132_839));
   MUX2_X1 i_132_0_121 (.A(\o_buffer[51] [6]), .B(i_mem_data[6]), .S(n_68), 
      .Z(n_132_838));
   MUX2_X1 i_132_0_122 (.A(\o_buffer[51] [5]), .B(i_mem_data[5]), .S(n_68), 
      .Z(n_132_837));
   MUX2_X1 i_132_0_123 (.A(\o_buffer[51] [4]), .B(i_mem_data[4]), .S(n_68), 
      .Z(n_132_836));
   MUX2_X1 i_132_0_124 (.A(\o_buffer[51] [3]), .B(i_mem_data[3]), .S(n_68), 
      .Z(n_132_835));
   MUX2_X1 i_132_0_125 (.A(\o_buffer[51] [2]), .B(i_mem_data[2]), .S(n_68), 
      .Z(n_132_834));
   MUX2_X1 i_132_0_126 (.A(\o_buffer[51] [1]), .B(i_mem_data[1]), .S(n_68), 
      .Z(n_132_833));
   MUX2_X1 i_132_0_127 (.A(\o_buffer[51] [0]), .B(i_mem_data[0]), .S(n_68), 
      .Z(n_132_832));
   MUX2_X1 i_132_0_128 (.A(\o_buffer[50] [15]), .B(i_mem_data[15]), .S(n_69), 
      .Z(n_132_831));
   MUX2_X1 i_132_0_129 (.A(\o_buffer[50] [14]), .B(i_mem_data[14]), .S(n_69), 
      .Z(n_132_830));
   MUX2_X1 i_132_0_130 (.A(\o_buffer[50] [13]), .B(i_mem_data[13]), .S(n_69), 
      .Z(n_132_829));
   MUX2_X1 i_132_0_131 (.A(\o_buffer[50] [12]), .B(i_mem_data[12]), .S(n_69), 
      .Z(n_132_828));
   MUX2_X1 i_132_0_132 (.A(\o_buffer[50] [11]), .B(i_mem_data[11]), .S(n_69), 
      .Z(n_132_827));
   MUX2_X1 i_132_0_133 (.A(\o_buffer[50] [10]), .B(i_mem_data[10]), .S(n_69), 
      .Z(n_132_826));
   MUX2_X1 i_132_0_134 (.A(\o_buffer[50] [9]), .B(i_mem_data[9]), .S(n_69), 
      .Z(n_132_825));
   MUX2_X1 i_132_0_135 (.A(\o_buffer[50] [8]), .B(i_mem_data[8]), .S(n_69), 
      .Z(n_132_824));
   MUX2_X1 i_132_0_136 (.A(\o_buffer[50] [7]), .B(i_mem_data[7]), .S(n_69), 
      .Z(n_132_823));
   MUX2_X1 i_132_0_137 (.A(\o_buffer[50] [6]), .B(i_mem_data[6]), .S(n_69), 
      .Z(n_132_822));
   MUX2_X1 i_132_0_138 (.A(\o_buffer[50] [5]), .B(i_mem_data[5]), .S(n_69), 
      .Z(n_132_821));
   MUX2_X1 i_132_0_139 (.A(\o_buffer[50] [4]), .B(i_mem_data[4]), .S(n_69), 
      .Z(n_132_820));
   MUX2_X1 i_132_0_140 (.A(\o_buffer[50] [3]), .B(i_mem_data[3]), .S(n_69), 
      .Z(n_132_819));
   MUX2_X1 i_132_0_141 (.A(\o_buffer[50] [2]), .B(i_mem_data[2]), .S(n_69), 
      .Z(n_132_818));
   MUX2_X1 i_132_0_142 (.A(\o_buffer[50] [1]), .B(i_mem_data[1]), .S(n_69), 
      .Z(n_132_817));
   MUX2_X1 i_132_0_143 (.A(\o_buffer[50] [0]), .B(i_mem_data[0]), .S(n_69), 
      .Z(n_132_816));
   MUX2_X1 i_132_0_144 (.A(\o_buffer[49] [15]), .B(i_mem_data[15]), .S(n_70), 
      .Z(n_132_815));
   MUX2_X1 i_132_0_145 (.A(\o_buffer[49] [14]), .B(i_mem_data[14]), .S(n_70), 
      .Z(n_132_814));
   MUX2_X1 i_132_0_146 (.A(\o_buffer[49] [13]), .B(i_mem_data[13]), .S(n_70), 
      .Z(n_132_813));
   MUX2_X1 i_132_0_147 (.A(\o_buffer[49] [12]), .B(i_mem_data[12]), .S(n_70), 
      .Z(n_132_812));
   MUX2_X1 i_132_0_148 (.A(\o_buffer[49] [11]), .B(i_mem_data[11]), .S(n_70), 
      .Z(n_132_811));
   MUX2_X1 i_132_0_149 (.A(\o_buffer[49] [10]), .B(i_mem_data[10]), .S(n_70), 
      .Z(n_132_810));
   MUX2_X1 i_132_0_150 (.A(\o_buffer[49] [9]), .B(i_mem_data[9]), .S(n_70), 
      .Z(n_132_809));
   MUX2_X1 i_132_0_151 (.A(\o_buffer[49] [8]), .B(i_mem_data[8]), .S(n_70), 
      .Z(n_132_808));
   MUX2_X1 i_132_0_152 (.A(\o_buffer[49] [7]), .B(i_mem_data[7]), .S(n_70), 
      .Z(n_132_807));
   MUX2_X1 i_132_0_153 (.A(\o_buffer[49] [6]), .B(i_mem_data[6]), .S(n_70), 
      .Z(n_132_806));
   MUX2_X1 i_132_0_154 (.A(\o_buffer[49] [5]), .B(i_mem_data[5]), .S(n_70), 
      .Z(n_132_805));
   MUX2_X1 i_132_0_155 (.A(\o_buffer[49] [4]), .B(i_mem_data[4]), .S(n_70), 
      .Z(n_132_804));
   MUX2_X1 i_132_0_156 (.A(\o_buffer[49] [3]), .B(i_mem_data[3]), .S(n_70), 
      .Z(n_132_803));
   MUX2_X1 i_132_0_157 (.A(\o_buffer[49] [2]), .B(i_mem_data[2]), .S(n_70), 
      .Z(n_132_802));
   MUX2_X1 i_132_0_158 (.A(\o_buffer[49] [1]), .B(i_mem_data[1]), .S(n_70), 
      .Z(n_132_801));
   MUX2_X1 i_132_0_159 (.A(\o_buffer[49] [0]), .B(i_mem_data[0]), .S(n_70), 
      .Z(n_132_800));
   MUX2_X1 i_132_0_160 (.A(\o_buffer[48] [15]), .B(i_mem_data[15]), .S(n_71), 
      .Z(n_132_799));
   MUX2_X1 i_132_0_161 (.A(\o_buffer[48] [14]), .B(i_mem_data[14]), .S(n_71), 
      .Z(n_132_798));
   MUX2_X1 i_132_0_162 (.A(\o_buffer[48] [13]), .B(i_mem_data[13]), .S(n_71), 
      .Z(n_132_797));
   MUX2_X1 i_132_0_163 (.A(\o_buffer[48] [12]), .B(i_mem_data[12]), .S(n_71), 
      .Z(n_132_796));
   MUX2_X1 i_132_0_164 (.A(\o_buffer[48] [11]), .B(i_mem_data[11]), .S(n_71), 
      .Z(n_132_795));
   MUX2_X1 i_132_0_165 (.A(\o_buffer[48] [10]), .B(i_mem_data[10]), .S(n_71), 
      .Z(n_132_794));
   MUX2_X1 i_132_0_166 (.A(\o_buffer[48] [9]), .B(i_mem_data[9]), .S(n_71), 
      .Z(n_132_793));
   MUX2_X1 i_132_0_167 (.A(\o_buffer[48] [8]), .B(i_mem_data[8]), .S(n_71), 
      .Z(n_132_792));
   MUX2_X1 i_132_0_168 (.A(\o_buffer[48] [7]), .B(i_mem_data[7]), .S(n_71), 
      .Z(n_132_791));
   MUX2_X1 i_132_0_169 (.A(\o_buffer[48] [6]), .B(i_mem_data[6]), .S(n_71), 
      .Z(n_132_790));
   MUX2_X1 i_132_0_170 (.A(\o_buffer[48] [5]), .B(i_mem_data[5]), .S(n_71), 
      .Z(n_132_789));
   MUX2_X1 i_132_0_171 (.A(\o_buffer[48] [4]), .B(i_mem_data[4]), .S(n_71), 
      .Z(n_132_788));
   MUX2_X1 i_132_0_172 (.A(\o_buffer[48] [3]), .B(i_mem_data[3]), .S(n_71), 
      .Z(n_132_787));
   MUX2_X1 i_132_0_173 (.A(\o_buffer[48] [2]), .B(i_mem_data[2]), .S(n_71), 
      .Z(n_132_786));
   MUX2_X1 i_132_0_174 (.A(\o_buffer[48] [1]), .B(i_mem_data[1]), .S(n_71), 
      .Z(n_132_785));
   MUX2_X1 i_132_0_175 (.A(\o_buffer[48] [0]), .B(i_mem_data[0]), .S(n_71), 
      .Z(n_132_784));
   MUX2_X1 i_132_0_176 (.A(\o_buffer[47] [15]), .B(i_mem_data[15]), .S(n_72), 
      .Z(n_132_783));
   MUX2_X1 i_132_0_177 (.A(\o_buffer[47] [14]), .B(i_mem_data[14]), .S(n_72), 
      .Z(n_132_782));
   MUX2_X1 i_132_0_178 (.A(\o_buffer[47] [13]), .B(i_mem_data[13]), .S(n_72), 
      .Z(n_132_781));
   MUX2_X1 i_132_0_179 (.A(\o_buffer[47] [12]), .B(i_mem_data[12]), .S(n_72), 
      .Z(n_132_780));
   MUX2_X1 i_132_0_180 (.A(\o_buffer[47] [11]), .B(i_mem_data[11]), .S(n_72), 
      .Z(n_132_779));
   MUX2_X1 i_132_0_181 (.A(\o_buffer[47] [10]), .B(i_mem_data[10]), .S(n_72), 
      .Z(n_132_778));
   MUX2_X1 i_132_0_182 (.A(\o_buffer[47] [9]), .B(i_mem_data[9]), .S(n_72), 
      .Z(n_132_777));
   MUX2_X1 i_132_0_183 (.A(\o_buffer[47] [8]), .B(i_mem_data[8]), .S(n_72), 
      .Z(n_132_776));
   MUX2_X1 i_132_0_184 (.A(\o_buffer[47] [7]), .B(i_mem_data[7]), .S(n_72), 
      .Z(n_132_775));
   MUX2_X1 i_132_0_185 (.A(\o_buffer[47] [6]), .B(i_mem_data[6]), .S(n_72), 
      .Z(n_132_774));
   MUX2_X1 i_132_0_186 (.A(\o_buffer[47] [5]), .B(i_mem_data[5]), .S(n_72), 
      .Z(n_132_773));
   MUX2_X1 i_132_0_187 (.A(\o_buffer[47] [4]), .B(i_mem_data[4]), .S(n_72), 
      .Z(n_132_772));
   MUX2_X1 i_132_0_188 (.A(\o_buffer[47] [3]), .B(i_mem_data[3]), .S(n_72), 
      .Z(n_132_771));
   MUX2_X1 i_132_0_189 (.A(\o_buffer[47] [2]), .B(i_mem_data[2]), .S(n_72), 
      .Z(n_132_770));
   MUX2_X1 i_132_0_190 (.A(\o_buffer[47] [1]), .B(i_mem_data[1]), .S(n_72), 
      .Z(n_132_769));
   MUX2_X1 i_132_0_191 (.A(\o_buffer[47] [0]), .B(i_mem_data[0]), .S(n_72), 
      .Z(n_132_768));
   MUX2_X1 i_132_0_192 (.A(\o_buffer[46] [15]), .B(i_mem_data[15]), .S(n_73), 
      .Z(n_132_767));
   MUX2_X1 i_132_0_193 (.A(\o_buffer[46] [14]), .B(i_mem_data[14]), .S(n_73), 
      .Z(n_132_766));
   MUX2_X1 i_132_0_194 (.A(\o_buffer[46] [13]), .B(i_mem_data[13]), .S(n_73), 
      .Z(n_132_765));
   MUX2_X1 i_132_0_195 (.A(\o_buffer[46] [12]), .B(i_mem_data[12]), .S(n_73), 
      .Z(n_132_764));
   MUX2_X1 i_132_0_196 (.A(\o_buffer[46] [11]), .B(i_mem_data[11]), .S(n_73), 
      .Z(n_132_763));
   MUX2_X1 i_132_0_197 (.A(\o_buffer[46] [10]), .B(i_mem_data[10]), .S(n_73), 
      .Z(n_132_762));
   MUX2_X1 i_132_0_198 (.A(\o_buffer[46] [9]), .B(i_mem_data[9]), .S(n_73), 
      .Z(n_132_761));
   MUX2_X1 i_132_0_199 (.A(\o_buffer[46] [8]), .B(i_mem_data[8]), .S(n_73), 
      .Z(n_132_760));
   MUX2_X1 i_132_0_200 (.A(\o_buffer[46] [7]), .B(i_mem_data[7]), .S(n_73), 
      .Z(n_132_759));
   MUX2_X1 i_132_0_201 (.A(\o_buffer[46] [6]), .B(i_mem_data[6]), .S(n_73), 
      .Z(n_132_758));
   MUX2_X1 i_132_0_202 (.A(\o_buffer[46] [5]), .B(i_mem_data[5]), .S(n_73), 
      .Z(n_132_757));
   MUX2_X1 i_132_0_203 (.A(\o_buffer[46] [4]), .B(i_mem_data[4]), .S(n_73), 
      .Z(n_132_756));
   MUX2_X1 i_132_0_204 (.A(\o_buffer[46] [3]), .B(i_mem_data[3]), .S(n_73), 
      .Z(n_132_755));
   MUX2_X1 i_132_0_205 (.A(\o_buffer[46] [2]), .B(i_mem_data[2]), .S(n_73), 
      .Z(n_132_754));
   MUX2_X1 i_132_0_206 (.A(\o_buffer[46] [1]), .B(i_mem_data[1]), .S(n_73), 
      .Z(n_132_753));
   MUX2_X1 i_132_0_207 (.A(\o_buffer[46] [0]), .B(i_mem_data[0]), .S(n_73), 
      .Z(n_132_752));
   MUX2_X1 i_132_0_208 (.A(\o_buffer[45] [15]), .B(i_mem_data[15]), .S(n_74), 
      .Z(n_132_751));
   MUX2_X1 i_132_0_209 (.A(\o_buffer[45] [14]), .B(i_mem_data[14]), .S(n_74), 
      .Z(n_132_750));
   MUX2_X1 i_132_0_210 (.A(\o_buffer[45] [13]), .B(i_mem_data[13]), .S(n_74), 
      .Z(n_132_749));
   MUX2_X1 i_132_0_211 (.A(\o_buffer[45] [12]), .B(i_mem_data[12]), .S(n_74), 
      .Z(n_132_748));
   MUX2_X1 i_132_0_212 (.A(\o_buffer[45] [11]), .B(i_mem_data[11]), .S(n_74), 
      .Z(n_132_747));
   MUX2_X1 i_132_0_213 (.A(\o_buffer[45] [10]), .B(i_mem_data[10]), .S(n_74), 
      .Z(n_132_746));
   MUX2_X1 i_132_0_214 (.A(\o_buffer[45] [9]), .B(i_mem_data[9]), .S(n_74), 
      .Z(n_132_745));
   MUX2_X1 i_132_0_215 (.A(\o_buffer[45] [8]), .B(i_mem_data[8]), .S(n_74), 
      .Z(n_132_744));
   MUX2_X1 i_132_0_216 (.A(\o_buffer[45] [7]), .B(i_mem_data[7]), .S(n_74), 
      .Z(n_132_743));
   MUX2_X1 i_132_0_217 (.A(\o_buffer[45] [6]), .B(i_mem_data[6]), .S(n_74), 
      .Z(n_132_742));
   MUX2_X1 i_132_0_218 (.A(\o_buffer[45] [5]), .B(i_mem_data[5]), .S(n_74), 
      .Z(n_132_741));
   MUX2_X1 i_132_0_219 (.A(\o_buffer[45] [4]), .B(i_mem_data[4]), .S(n_74), 
      .Z(n_132_740));
   MUX2_X1 i_132_0_220 (.A(\o_buffer[45] [3]), .B(i_mem_data[3]), .S(n_74), 
      .Z(n_132_739));
   MUX2_X1 i_132_0_221 (.A(\o_buffer[45] [2]), .B(i_mem_data[2]), .S(n_74), 
      .Z(n_132_738));
   MUX2_X1 i_132_0_222 (.A(\o_buffer[45] [1]), .B(i_mem_data[1]), .S(n_74), 
      .Z(n_132_737));
   MUX2_X1 i_132_0_223 (.A(\o_buffer[45] [0]), .B(i_mem_data[0]), .S(n_74), 
      .Z(n_132_736));
   MUX2_X1 i_132_0_224 (.A(\o_buffer[44] [15]), .B(i_mem_data[15]), .S(n_75), 
      .Z(n_132_735));
   MUX2_X1 i_132_0_225 (.A(\o_buffer[44] [14]), .B(i_mem_data[14]), .S(n_75), 
      .Z(n_132_734));
   MUX2_X1 i_132_0_226 (.A(\o_buffer[44] [13]), .B(i_mem_data[13]), .S(n_75), 
      .Z(n_132_733));
   MUX2_X1 i_132_0_227 (.A(\o_buffer[44] [12]), .B(i_mem_data[12]), .S(n_75), 
      .Z(n_132_732));
   MUX2_X1 i_132_0_228 (.A(\o_buffer[44] [11]), .B(i_mem_data[11]), .S(n_75), 
      .Z(n_132_731));
   MUX2_X1 i_132_0_229 (.A(\o_buffer[44] [10]), .B(i_mem_data[10]), .S(n_75), 
      .Z(n_132_730));
   MUX2_X1 i_132_0_230 (.A(\o_buffer[44] [9]), .B(i_mem_data[9]), .S(n_75), 
      .Z(n_132_729));
   MUX2_X1 i_132_0_231 (.A(\o_buffer[44] [8]), .B(i_mem_data[8]), .S(n_75), 
      .Z(n_132_728));
   MUX2_X1 i_132_0_232 (.A(\o_buffer[44] [7]), .B(i_mem_data[7]), .S(n_75), 
      .Z(n_132_727));
   MUX2_X1 i_132_0_233 (.A(\o_buffer[44] [6]), .B(i_mem_data[6]), .S(n_75), 
      .Z(n_132_726));
   MUX2_X1 i_132_0_234 (.A(\o_buffer[44] [5]), .B(i_mem_data[5]), .S(n_75), 
      .Z(n_132_725));
   MUX2_X1 i_132_0_235 (.A(\o_buffer[44] [4]), .B(i_mem_data[4]), .S(n_75), 
      .Z(n_132_724));
   MUX2_X1 i_132_0_236 (.A(\o_buffer[44] [3]), .B(i_mem_data[3]), .S(n_75), 
      .Z(n_132_723));
   MUX2_X1 i_132_0_237 (.A(\o_buffer[44] [2]), .B(i_mem_data[2]), .S(n_75), 
      .Z(n_132_722));
   MUX2_X1 i_132_0_238 (.A(\o_buffer[44] [1]), .B(i_mem_data[1]), .S(n_75), 
      .Z(n_132_721));
   MUX2_X1 i_132_0_239 (.A(\o_buffer[44] [0]), .B(i_mem_data[0]), .S(n_75), 
      .Z(n_132_720));
   MUX2_X1 i_132_0_240 (.A(\o_buffer[43] [15]), .B(i_mem_data[15]), .S(n_76), 
      .Z(n_132_719));
   MUX2_X1 i_132_0_241 (.A(\o_buffer[43] [14]), .B(i_mem_data[14]), .S(n_76), 
      .Z(n_132_718));
   MUX2_X1 i_132_0_242 (.A(\o_buffer[43] [13]), .B(i_mem_data[13]), .S(n_76), 
      .Z(n_132_717));
   MUX2_X1 i_132_0_243 (.A(\o_buffer[43] [12]), .B(i_mem_data[12]), .S(n_76), 
      .Z(n_132_716));
   MUX2_X1 i_132_0_244 (.A(\o_buffer[43] [11]), .B(i_mem_data[11]), .S(n_76), 
      .Z(n_132_715));
   MUX2_X1 i_132_0_245 (.A(\o_buffer[43] [10]), .B(i_mem_data[10]), .S(n_76), 
      .Z(n_132_714));
   MUX2_X1 i_132_0_246 (.A(\o_buffer[43] [9]), .B(i_mem_data[9]), .S(n_76), 
      .Z(n_132_713));
   MUX2_X1 i_132_0_247 (.A(\o_buffer[43] [8]), .B(i_mem_data[8]), .S(n_76), 
      .Z(n_132_712));
   MUX2_X1 i_132_0_248 (.A(\o_buffer[43] [7]), .B(i_mem_data[7]), .S(n_76), 
      .Z(n_132_711));
   MUX2_X1 i_132_0_249 (.A(\o_buffer[43] [6]), .B(i_mem_data[6]), .S(n_76), 
      .Z(n_132_710));
   MUX2_X1 i_132_0_250 (.A(\o_buffer[43] [5]), .B(i_mem_data[5]), .S(n_76), 
      .Z(n_132_709));
   MUX2_X1 i_132_0_251 (.A(\o_buffer[43] [4]), .B(i_mem_data[4]), .S(n_76), 
      .Z(n_132_708));
   MUX2_X1 i_132_0_252 (.A(\o_buffer[43] [3]), .B(i_mem_data[3]), .S(n_76), 
      .Z(n_132_707));
   MUX2_X1 i_132_0_253 (.A(\o_buffer[43] [2]), .B(i_mem_data[2]), .S(n_76), 
      .Z(n_132_706));
   MUX2_X1 i_132_0_254 (.A(\o_buffer[43] [1]), .B(i_mem_data[1]), .S(n_76), 
      .Z(n_132_705));
   MUX2_X1 i_132_0_255 (.A(\o_buffer[43] [0]), .B(i_mem_data[0]), .S(n_76), 
      .Z(n_132_704));
   MUX2_X1 i_132_0_256 (.A(\o_buffer[42] [15]), .B(i_mem_data[15]), .S(n_77), 
      .Z(n_132_703));
   MUX2_X1 i_132_0_257 (.A(\o_buffer[42] [14]), .B(i_mem_data[14]), .S(n_77), 
      .Z(n_132_702));
   MUX2_X1 i_132_0_258 (.A(\o_buffer[42] [13]), .B(i_mem_data[13]), .S(n_77), 
      .Z(n_132_701));
   MUX2_X1 i_132_0_259 (.A(\o_buffer[42] [12]), .B(i_mem_data[12]), .S(n_77), 
      .Z(n_132_700));
   MUX2_X1 i_132_0_260 (.A(\o_buffer[42] [11]), .B(i_mem_data[11]), .S(n_77), 
      .Z(n_132_699));
   MUX2_X1 i_132_0_261 (.A(\o_buffer[42] [10]), .B(i_mem_data[10]), .S(n_77), 
      .Z(n_132_698));
   MUX2_X1 i_132_0_262 (.A(\o_buffer[42] [9]), .B(i_mem_data[9]), .S(n_77), 
      .Z(n_132_697));
   MUX2_X1 i_132_0_263 (.A(\o_buffer[42] [8]), .B(i_mem_data[8]), .S(n_77), 
      .Z(n_132_696));
   MUX2_X1 i_132_0_264 (.A(\o_buffer[42] [7]), .B(i_mem_data[7]), .S(n_77), 
      .Z(n_132_695));
   MUX2_X1 i_132_0_265 (.A(\o_buffer[42] [6]), .B(i_mem_data[6]), .S(n_77), 
      .Z(n_132_694));
   MUX2_X1 i_132_0_266 (.A(\o_buffer[42] [5]), .B(i_mem_data[5]), .S(n_77), 
      .Z(n_132_693));
   MUX2_X1 i_132_0_267 (.A(\o_buffer[42] [4]), .B(i_mem_data[4]), .S(n_77), 
      .Z(n_132_692));
   MUX2_X1 i_132_0_268 (.A(\o_buffer[42] [3]), .B(i_mem_data[3]), .S(n_77), 
      .Z(n_132_691));
   MUX2_X1 i_132_0_269 (.A(\o_buffer[42] [2]), .B(i_mem_data[2]), .S(n_77), 
      .Z(n_132_690));
   MUX2_X1 i_132_0_270 (.A(\o_buffer[42] [1]), .B(i_mem_data[1]), .S(n_77), 
      .Z(n_132_689));
   MUX2_X1 i_132_0_271 (.A(\o_buffer[42] [0]), .B(i_mem_data[0]), .S(n_77), 
      .Z(n_132_688));
   MUX2_X1 i_132_0_272 (.A(\o_buffer[41] [15]), .B(i_mem_data[15]), .S(n_78), 
      .Z(n_132_687));
   MUX2_X1 i_132_0_273 (.A(\o_buffer[41] [14]), .B(i_mem_data[14]), .S(n_78), 
      .Z(n_132_686));
   MUX2_X1 i_132_0_274 (.A(\o_buffer[41] [13]), .B(i_mem_data[13]), .S(n_78), 
      .Z(n_132_685));
   MUX2_X1 i_132_0_275 (.A(\o_buffer[41] [12]), .B(i_mem_data[12]), .S(n_78), 
      .Z(n_132_684));
   MUX2_X1 i_132_0_276 (.A(\o_buffer[41] [11]), .B(i_mem_data[11]), .S(n_78), 
      .Z(n_132_683));
   MUX2_X1 i_132_0_277 (.A(\o_buffer[41] [10]), .B(i_mem_data[10]), .S(n_78), 
      .Z(n_132_682));
   MUX2_X1 i_132_0_278 (.A(\o_buffer[41] [9]), .B(i_mem_data[9]), .S(n_78), 
      .Z(n_132_681));
   MUX2_X1 i_132_0_279 (.A(\o_buffer[41] [8]), .B(i_mem_data[8]), .S(n_78), 
      .Z(n_132_680));
   MUX2_X1 i_132_0_280 (.A(\o_buffer[41] [7]), .B(i_mem_data[7]), .S(n_78), 
      .Z(n_132_679));
   MUX2_X1 i_132_0_281 (.A(\o_buffer[41] [6]), .B(i_mem_data[6]), .S(n_78), 
      .Z(n_132_678));
   MUX2_X1 i_132_0_282 (.A(\o_buffer[41] [5]), .B(i_mem_data[5]), .S(n_78), 
      .Z(n_132_677));
   MUX2_X1 i_132_0_283 (.A(\o_buffer[41] [4]), .B(i_mem_data[4]), .S(n_78), 
      .Z(n_132_676));
   MUX2_X1 i_132_0_284 (.A(\o_buffer[41] [3]), .B(i_mem_data[3]), .S(n_78), 
      .Z(n_132_675));
   MUX2_X1 i_132_0_285 (.A(\o_buffer[41] [2]), .B(i_mem_data[2]), .S(n_78), 
      .Z(n_132_674));
   MUX2_X1 i_132_0_286 (.A(\o_buffer[41] [1]), .B(i_mem_data[1]), .S(n_78), 
      .Z(n_132_673));
   MUX2_X1 i_132_0_287 (.A(\o_buffer[41] [0]), .B(i_mem_data[0]), .S(n_78), 
      .Z(n_132_672));
   MUX2_X1 i_132_0_288 (.A(\o_buffer[40] [15]), .B(i_mem_data[15]), .S(n_79), 
      .Z(n_132_671));
   MUX2_X1 i_132_0_289 (.A(\o_buffer[40] [14]), .B(i_mem_data[14]), .S(n_79), 
      .Z(n_132_670));
   MUX2_X1 i_132_0_290 (.A(\o_buffer[40] [13]), .B(i_mem_data[13]), .S(n_79), 
      .Z(n_132_669));
   MUX2_X1 i_132_0_291 (.A(\o_buffer[40] [12]), .B(i_mem_data[12]), .S(n_79), 
      .Z(n_132_668));
   MUX2_X1 i_132_0_292 (.A(\o_buffer[40] [11]), .B(i_mem_data[11]), .S(n_79), 
      .Z(n_132_667));
   MUX2_X1 i_132_0_293 (.A(\o_buffer[40] [10]), .B(i_mem_data[10]), .S(n_79), 
      .Z(n_132_666));
   MUX2_X1 i_132_0_294 (.A(\o_buffer[40] [9]), .B(i_mem_data[9]), .S(n_79), 
      .Z(n_132_665));
   MUX2_X1 i_132_0_295 (.A(\o_buffer[40] [8]), .B(i_mem_data[8]), .S(n_79), 
      .Z(n_132_664));
   MUX2_X1 i_132_0_296 (.A(\o_buffer[40] [7]), .B(i_mem_data[7]), .S(n_79), 
      .Z(n_132_663));
   MUX2_X1 i_132_0_297 (.A(\o_buffer[40] [6]), .B(i_mem_data[6]), .S(n_79), 
      .Z(n_132_662));
   MUX2_X1 i_132_0_298 (.A(\o_buffer[40] [5]), .B(i_mem_data[5]), .S(n_79), 
      .Z(n_132_661));
   MUX2_X1 i_132_0_299 (.A(\o_buffer[40] [4]), .B(i_mem_data[4]), .S(n_79), 
      .Z(n_132_660));
   MUX2_X1 i_132_0_300 (.A(\o_buffer[40] [3]), .B(i_mem_data[3]), .S(n_79), 
      .Z(n_132_659));
   MUX2_X1 i_132_0_301 (.A(\o_buffer[40] [2]), .B(i_mem_data[2]), .S(n_79), 
      .Z(n_132_658));
   MUX2_X1 i_132_0_302 (.A(\o_buffer[40] [1]), .B(i_mem_data[1]), .S(n_79), 
      .Z(n_132_657));
   MUX2_X1 i_132_0_303 (.A(\o_buffer[40] [0]), .B(i_mem_data[0]), .S(n_79), 
      .Z(n_132_656));
   MUX2_X1 i_132_0_304 (.A(\o_buffer[39] [15]), .B(i_mem_data[15]), .S(n_80), 
      .Z(n_132_655));
   MUX2_X1 i_132_0_305 (.A(\o_buffer[39] [14]), .B(i_mem_data[14]), .S(n_80), 
      .Z(n_132_654));
   MUX2_X1 i_132_0_306 (.A(\o_buffer[39] [13]), .B(i_mem_data[13]), .S(n_80), 
      .Z(n_132_653));
   MUX2_X1 i_132_0_307 (.A(\o_buffer[39] [12]), .B(i_mem_data[12]), .S(n_80), 
      .Z(n_132_652));
   MUX2_X1 i_132_0_308 (.A(\o_buffer[39] [11]), .B(i_mem_data[11]), .S(n_80), 
      .Z(n_132_651));
   MUX2_X1 i_132_0_309 (.A(\o_buffer[39] [10]), .B(i_mem_data[10]), .S(n_80), 
      .Z(n_132_650));
   MUX2_X1 i_132_0_310 (.A(\o_buffer[39] [9]), .B(i_mem_data[9]), .S(n_80), 
      .Z(n_132_649));
   MUX2_X1 i_132_0_311 (.A(\o_buffer[39] [8]), .B(i_mem_data[8]), .S(n_80), 
      .Z(n_132_648));
   MUX2_X1 i_132_0_312 (.A(\o_buffer[39] [7]), .B(i_mem_data[7]), .S(n_80), 
      .Z(n_132_647));
   MUX2_X1 i_132_0_313 (.A(\o_buffer[39] [6]), .B(i_mem_data[6]), .S(n_80), 
      .Z(n_132_646));
   MUX2_X1 i_132_0_314 (.A(\o_buffer[39] [5]), .B(i_mem_data[5]), .S(n_80), 
      .Z(n_132_645));
   MUX2_X1 i_132_0_315 (.A(\o_buffer[39] [4]), .B(i_mem_data[4]), .S(n_80), 
      .Z(n_132_644));
   MUX2_X1 i_132_0_316 (.A(\o_buffer[39] [3]), .B(i_mem_data[3]), .S(n_80), 
      .Z(n_132_643));
   MUX2_X1 i_132_0_317 (.A(\o_buffer[39] [2]), .B(i_mem_data[2]), .S(n_80), 
      .Z(n_132_642));
   MUX2_X1 i_132_0_318 (.A(\o_buffer[39] [1]), .B(i_mem_data[1]), .S(n_80), 
      .Z(n_132_641));
   MUX2_X1 i_132_0_319 (.A(\o_buffer[39] [0]), .B(i_mem_data[0]), .S(n_80), 
      .Z(n_132_640));
   MUX2_X1 i_132_0_320 (.A(\o_buffer[38] [15]), .B(i_mem_data[15]), .S(n_81), 
      .Z(n_132_639));
   MUX2_X1 i_132_0_321 (.A(\o_buffer[38] [14]), .B(i_mem_data[14]), .S(n_81), 
      .Z(n_132_638));
   MUX2_X1 i_132_0_322 (.A(\o_buffer[38] [13]), .B(i_mem_data[13]), .S(n_81), 
      .Z(n_132_637));
   MUX2_X1 i_132_0_323 (.A(\o_buffer[38] [12]), .B(i_mem_data[12]), .S(n_81), 
      .Z(n_132_636));
   MUX2_X1 i_132_0_324 (.A(\o_buffer[38] [11]), .B(i_mem_data[11]), .S(n_81), 
      .Z(n_132_635));
   MUX2_X1 i_132_0_325 (.A(\o_buffer[38] [10]), .B(i_mem_data[10]), .S(n_81), 
      .Z(n_132_634));
   MUX2_X1 i_132_0_326 (.A(\o_buffer[38] [9]), .B(i_mem_data[9]), .S(n_81), 
      .Z(n_132_633));
   MUX2_X1 i_132_0_327 (.A(\o_buffer[38] [8]), .B(i_mem_data[8]), .S(n_81), 
      .Z(n_132_632));
   MUX2_X1 i_132_0_328 (.A(\o_buffer[38] [7]), .B(i_mem_data[7]), .S(n_81), 
      .Z(n_132_631));
   MUX2_X1 i_132_0_329 (.A(\o_buffer[38] [6]), .B(i_mem_data[6]), .S(n_81), 
      .Z(n_132_630));
   MUX2_X1 i_132_0_330 (.A(\o_buffer[38] [5]), .B(i_mem_data[5]), .S(n_81), 
      .Z(n_132_629));
   MUX2_X1 i_132_0_331 (.A(\o_buffer[38] [4]), .B(i_mem_data[4]), .S(n_81), 
      .Z(n_132_628));
   MUX2_X1 i_132_0_332 (.A(\o_buffer[38] [3]), .B(i_mem_data[3]), .S(n_81), 
      .Z(n_132_627));
   MUX2_X1 i_132_0_333 (.A(\o_buffer[38] [2]), .B(i_mem_data[2]), .S(n_81), 
      .Z(n_132_626));
   MUX2_X1 i_132_0_334 (.A(\o_buffer[38] [1]), .B(i_mem_data[1]), .S(n_81), 
      .Z(n_132_625));
   MUX2_X1 i_132_0_335 (.A(\o_buffer[38] [0]), .B(i_mem_data[0]), .S(n_81), 
      .Z(n_132_624));
   MUX2_X1 i_132_0_336 (.A(\o_buffer[37] [15]), .B(i_mem_data[15]), .S(n_82), 
      .Z(n_132_623));
   MUX2_X1 i_132_0_337 (.A(\o_buffer[37] [14]), .B(i_mem_data[14]), .S(n_82), 
      .Z(n_132_622));
   MUX2_X1 i_132_0_338 (.A(\o_buffer[37] [13]), .B(i_mem_data[13]), .S(n_82), 
      .Z(n_132_621));
   MUX2_X1 i_132_0_339 (.A(\o_buffer[37] [12]), .B(i_mem_data[12]), .S(n_82), 
      .Z(n_132_620));
   MUX2_X1 i_132_0_340 (.A(\o_buffer[37] [11]), .B(i_mem_data[11]), .S(n_82), 
      .Z(n_132_619));
   MUX2_X1 i_132_0_341 (.A(\o_buffer[37] [10]), .B(i_mem_data[10]), .S(n_82), 
      .Z(n_132_618));
   MUX2_X1 i_132_0_342 (.A(\o_buffer[37] [9]), .B(i_mem_data[9]), .S(n_82), 
      .Z(n_132_617));
   MUX2_X1 i_132_0_343 (.A(\o_buffer[37] [8]), .B(i_mem_data[8]), .S(n_82), 
      .Z(n_132_616));
   MUX2_X1 i_132_0_344 (.A(\o_buffer[37] [7]), .B(i_mem_data[7]), .S(n_82), 
      .Z(n_132_615));
   MUX2_X1 i_132_0_345 (.A(\o_buffer[37] [6]), .B(i_mem_data[6]), .S(n_82), 
      .Z(n_132_614));
   MUX2_X1 i_132_0_346 (.A(\o_buffer[37] [5]), .B(i_mem_data[5]), .S(n_82), 
      .Z(n_132_613));
   MUX2_X1 i_132_0_347 (.A(\o_buffer[37] [4]), .B(i_mem_data[4]), .S(n_82), 
      .Z(n_132_612));
   MUX2_X1 i_132_0_348 (.A(\o_buffer[37] [3]), .B(i_mem_data[3]), .S(n_82), 
      .Z(n_132_611));
   MUX2_X1 i_132_0_349 (.A(\o_buffer[37] [2]), .B(i_mem_data[2]), .S(n_82), 
      .Z(n_132_610));
   MUX2_X1 i_132_0_350 (.A(\o_buffer[37] [1]), .B(i_mem_data[1]), .S(n_82), 
      .Z(n_132_609));
   MUX2_X1 i_132_0_351 (.A(\o_buffer[37] [0]), .B(i_mem_data[0]), .S(n_82), 
      .Z(n_132_608));
   MUX2_X1 i_132_0_352 (.A(\o_buffer[36] [15]), .B(i_mem_data[15]), .S(n_83), 
      .Z(n_132_607));
   MUX2_X1 i_132_0_353 (.A(\o_buffer[36] [14]), .B(i_mem_data[14]), .S(n_83), 
      .Z(n_132_606));
   MUX2_X1 i_132_0_354 (.A(\o_buffer[36] [13]), .B(i_mem_data[13]), .S(n_83), 
      .Z(n_132_605));
   MUX2_X1 i_132_0_355 (.A(\o_buffer[36] [12]), .B(i_mem_data[12]), .S(n_83), 
      .Z(n_132_604));
   MUX2_X1 i_132_0_356 (.A(\o_buffer[36] [11]), .B(i_mem_data[11]), .S(n_83), 
      .Z(n_132_603));
   MUX2_X1 i_132_0_357 (.A(\o_buffer[36] [10]), .B(i_mem_data[10]), .S(n_83), 
      .Z(n_132_602));
   MUX2_X1 i_132_0_358 (.A(\o_buffer[36] [9]), .B(i_mem_data[9]), .S(n_83), 
      .Z(n_132_601));
   MUX2_X1 i_132_0_359 (.A(\o_buffer[36] [8]), .B(i_mem_data[8]), .S(n_83), 
      .Z(n_132_600));
   MUX2_X1 i_132_0_360 (.A(\o_buffer[36] [7]), .B(i_mem_data[7]), .S(n_83), 
      .Z(n_132_599));
   MUX2_X1 i_132_0_361 (.A(\o_buffer[36] [6]), .B(i_mem_data[6]), .S(n_83), 
      .Z(n_132_598));
   MUX2_X1 i_132_0_362 (.A(\o_buffer[36] [5]), .B(i_mem_data[5]), .S(n_83), 
      .Z(n_132_597));
   MUX2_X1 i_132_0_363 (.A(\o_buffer[36] [4]), .B(i_mem_data[4]), .S(n_83), 
      .Z(n_132_596));
   MUX2_X1 i_132_0_364 (.A(\o_buffer[36] [3]), .B(i_mem_data[3]), .S(n_83), 
      .Z(n_132_595));
   MUX2_X1 i_132_0_365 (.A(\o_buffer[36] [2]), .B(i_mem_data[2]), .S(n_83), 
      .Z(n_132_594));
   MUX2_X1 i_132_0_366 (.A(\o_buffer[36] [1]), .B(i_mem_data[1]), .S(n_83), 
      .Z(n_132_593));
   MUX2_X1 i_132_0_367 (.A(\o_buffer[36] [0]), .B(i_mem_data[0]), .S(n_83), 
      .Z(n_132_592));
   MUX2_X1 i_132_0_368 (.A(\o_buffer[35] [15]), .B(i_mem_data[15]), .S(n_84), 
      .Z(n_132_591));
   MUX2_X1 i_132_0_369 (.A(\o_buffer[35] [14]), .B(i_mem_data[14]), .S(n_84), 
      .Z(n_132_590));
   MUX2_X1 i_132_0_370 (.A(\o_buffer[35] [13]), .B(i_mem_data[13]), .S(n_84), 
      .Z(n_132_589));
   MUX2_X1 i_132_0_371 (.A(\o_buffer[35] [12]), .B(i_mem_data[12]), .S(n_84), 
      .Z(n_132_588));
   MUX2_X1 i_132_0_372 (.A(\o_buffer[35] [11]), .B(i_mem_data[11]), .S(n_84), 
      .Z(n_132_587));
   MUX2_X1 i_132_0_373 (.A(\o_buffer[35] [10]), .B(i_mem_data[10]), .S(n_84), 
      .Z(n_132_586));
   MUX2_X1 i_132_0_374 (.A(\o_buffer[35] [9]), .B(i_mem_data[9]), .S(n_84), 
      .Z(n_132_585));
   MUX2_X1 i_132_0_375 (.A(\o_buffer[35] [8]), .B(i_mem_data[8]), .S(n_84), 
      .Z(n_132_584));
   MUX2_X1 i_132_0_376 (.A(\o_buffer[35] [7]), .B(i_mem_data[7]), .S(n_84), 
      .Z(n_132_583));
   MUX2_X1 i_132_0_377 (.A(\o_buffer[35] [6]), .B(i_mem_data[6]), .S(n_84), 
      .Z(n_132_582));
   MUX2_X1 i_132_0_378 (.A(\o_buffer[35] [5]), .B(i_mem_data[5]), .S(n_84), 
      .Z(n_132_581));
   MUX2_X1 i_132_0_379 (.A(\o_buffer[35] [4]), .B(i_mem_data[4]), .S(n_84), 
      .Z(n_132_580));
   MUX2_X1 i_132_0_380 (.A(\o_buffer[35] [3]), .B(i_mem_data[3]), .S(n_84), 
      .Z(n_132_579));
   MUX2_X1 i_132_0_381 (.A(\o_buffer[35] [2]), .B(i_mem_data[2]), .S(n_84), 
      .Z(n_132_578));
   MUX2_X1 i_132_0_382 (.A(\o_buffer[35] [1]), .B(i_mem_data[1]), .S(n_84), 
      .Z(n_132_577));
   MUX2_X1 i_132_0_383 (.A(\o_buffer[35] [0]), .B(i_mem_data[0]), .S(n_84), 
      .Z(n_132_576));
   MUX2_X1 i_132_0_384 (.A(\o_buffer[34] [15]), .B(i_mem_data[15]), .S(n_85), 
      .Z(n_132_575));
   MUX2_X1 i_132_0_385 (.A(\o_buffer[34] [14]), .B(i_mem_data[14]), .S(n_85), 
      .Z(n_132_574));
   MUX2_X1 i_132_0_386 (.A(\o_buffer[34] [13]), .B(i_mem_data[13]), .S(n_85), 
      .Z(n_132_573));
   MUX2_X1 i_132_0_387 (.A(\o_buffer[34] [12]), .B(i_mem_data[12]), .S(n_85), 
      .Z(n_132_572));
   MUX2_X1 i_132_0_388 (.A(\o_buffer[34] [11]), .B(i_mem_data[11]), .S(n_85), 
      .Z(n_132_571));
   MUX2_X1 i_132_0_389 (.A(\o_buffer[34] [10]), .B(i_mem_data[10]), .S(n_85), 
      .Z(n_132_570));
   MUX2_X1 i_132_0_390 (.A(\o_buffer[34] [9]), .B(i_mem_data[9]), .S(n_85), 
      .Z(n_132_569));
   MUX2_X1 i_132_0_391 (.A(\o_buffer[34] [8]), .B(i_mem_data[8]), .S(n_85), 
      .Z(n_132_568));
   MUX2_X1 i_132_0_392 (.A(\o_buffer[34] [7]), .B(i_mem_data[7]), .S(n_85), 
      .Z(n_132_567));
   MUX2_X1 i_132_0_393 (.A(\o_buffer[34] [6]), .B(i_mem_data[6]), .S(n_85), 
      .Z(n_132_566));
   MUX2_X1 i_132_0_394 (.A(\o_buffer[34] [5]), .B(i_mem_data[5]), .S(n_85), 
      .Z(n_132_565));
   MUX2_X1 i_132_0_395 (.A(\o_buffer[34] [4]), .B(i_mem_data[4]), .S(n_85), 
      .Z(n_132_564));
   MUX2_X1 i_132_0_396 (.A(\o_buffer[34] [3]), .B(i_mem_data[3]), .S(n_85), 
      .Z(n_132_563));
   MUX2_X1 i_132_0_397 (.A(\o_buffer[34] [2]), .B(i_mem_data[2]), .S(n_85), 
      .Z(n_132_562));
   MUX2_X1 i_132_0_398 (.A(\o_buffer[34] [1]), .B(i_mem_data[1]), .S(n_85), 
      .Z(n_132_561));
   MUX2_X1 i_132_0_399 (.A(\o_buffer[34] [0]), .B(i_mem_data[0]), .S(n_85), 
      .Z(n_132_560));
   MUX2_X1 i_132_0_400 (.A(\o_buffer[33] [15]), .B(i_mem_data[15]), .S(n_86), 
      .Z(n_132_559));
   MUX2_X1 i_132_0_401 (.A(\o_buffer[33] [14]), .B(i_mem_data[14]), .S(n_86), 
      .Z(n_132_558));
   MUX2_X1 i_132_0_402 (.A(\o_buffer[33] [13]), .B(i_mem_data[13]), .S(n_86), 
      .Z(n_132_557));
   MUX2_X1 i_132_0_403 (.A(\o_buffer[33] [12]), .B(i_mem_data[12]), .S(n_86), 
      .Z(n_132_556));
   MUX2_X1 i_132_0_404 (.A(\o_buffer[33] [11]), .B(i_mem_data[11]), .S(n_86), 
      .Z(n_132_555));
   MUX2_X1 i_132_0_405 (.A(\o_buffer[33] [10]), .B(i_mem_data[10]), .S(n_86), 
      .Z(n_132_554));
   MUX2_X1 i_132_0_406 (.A(\o_buffer[33] [9]), .B(i_mem_data[9]), .S(n_86), 
      .Z(n_132_553));
   MUX2_X1 i_132_0_407 (.A(\o_buffer[33] [8]), .B(i_mem_data[8]), .S(n_86), 
      .Z(n_132_552));
   MUX2_X1 i_132_0_408 (.A(\o_buffer[33] [7]), .B(i_mem_data[7]), .S(n_86), 
      .Z(n_132_551));
   MUX2_X1 i_132_0_409 (.A(\o_buffer[33] [6]), .B(i_mem_data[6]), .S(n_86), 
      .Z(n_132_550));
   MUX2_X1 i_132_0_410 (.A(\o_buffer[33] [5]), .B(i_mem_data[5]), .S(n_86), 
      .Z(n_132_549));
   MUX2_X1 i_132_0_411 (.A(\o_buffer[33] [4]), .B(i_mem_data[4]), .S(n_86), 
      .Z(n_132_548));
   MUX2_X1 i_132_0_412 (.A(\o_buffer[33] [3]), .B(i_mem_data[3]), .S(n_86), 
      .Z(n_132_547));
   MUX2_X1 i_132_0_413 (.A(\o_buffer[33] [2]), .B(i_mem_data[2]), .S(n_86), 
      .Z(n_132_546));
   MUX2_X1 i_132_0_414 (.A(\o_buffer[33] [1]), .B(i_mem_data[1]), .S(n_86), 
      .Z(n_132_545));
   MUX2_X1 i_132_0_415 (.A(\o_buffer[33] [0]), .B(i_mem_data[0]), .S(n_86), 
      .Z(n_132_544));
   MUX2_X1 i_132_0_416 (.A(\o_buffer[32] [15]), .B(i_mem_data[15]), .S(n_87), 
      .Z(n_132_543));
   MUX2_X1 i_132_0_417 (.A(\o_buffer[32] [14]), .B(i_mem_data[14]), .S(n_87), 
      .Z(n_132_542));
   MUX2_X1 i_132_0_418 (.A(\o_buffer[32] [13]), .B(i_mem_data[13]), .S(n_87), 
      .Z(n_132_541));
   MUX2_X1 i_132_0_419 (.A(\o_buffer[32] [12]), .B(i_mem_data[12]), .S(n_87), 
      .Z(n_132_540));
   MUX2_X1 i_132_0_420 (.A(\o_buffer[32] [11]), .B(i_mem_data[11]), .S(n_87), 
      .Z(n_132_539));
   MUX2_X1 i_132_0_421 (.A(\o_buffer[32] [10]), .B(i_mem_data[10]), .S(n_87), 
      .Z(n_132_538));
   MUX2_X1 i_132_0_422 (.A(\o_buffer[32] [9]), .B(i_mem_data[9]), .S(n_87), 
      .Z(n_132_537));
   MUX2_X1 i_132_0_423 (.A(\o_buffer[32] [8]), .B(i_mem_data[8]), .S(n_87), 
      .Z(n_132_536));
   MUX2_X1 i_132_0_424 (.A(\o_buffer[32] [7]), .B(i_mem_data[7]), .S(n_87), 
      .Z(n_132_535));
   MUX2_X1 i_132_0_425 (.A(\o_buffer[32] [6]), .B(i_mem_data[6]), .S(n_87), 
      .Z(n_132_534));
   MUX2_X1 i_132_0_426 (.A(\o_buffer[32] [5]), .B(i_mem_data[5]), .S(n_87), 
      .Z(n_132_533));
   MUX2_X1 i_132_0_427 (.A(\o_buffer[32] [4]), .B(i_mem_data[4]), .S(n_87), 
      .Z(n_132_532));
   MUX2_X1 i_132_0_428 (.A(\o_buffer[32] [3]), .B(i_mem_data[3]), .S(n_87), 
      .Z(n_132_531));
   MUX2_X1 i_132_0_429 (.A(\o_buffer[32] [2]), .B(i_mem_data[2]), .S(n_87), 
      .Z(n_132_530));
   MUX2_X1 i_132_0_430 (.A(\o_buffer[32] [1]), .B(i_mem_data[1]), .S(n_87), 
      .Z(n_132_529));
   MUX2_X1 i_132_0_431 (.A(\o_buffer[32] [0]), .B(i_mem_data[0]), .S(n_87), 
      .Z(n_132_528));
   MUX2_X1 i_132_0_432 (.A(\o_buffer[31] [15]), .B(i_mem_data[15]), .S(n_88), 
      .Z(n_132_527));
   MUX2_X1 i_132_0_433 (.A(\o_buffer[31] [14]), .B(i_mem_data[14]), .S(n_88), 
      .Z(n_132_526));
   MUX2_X1 i_132_0_434 (.A(\o_buffer[31] [13]), .B(i_mem_data[13]), .S(n_88), 
      .Z(n_132_525));
   MUX2_X1 i_132_0_435 (.A(\o_buffer[31] [12]), .B(i_mem_data[12]), .S(n_88), 
      .Z(n_132_524));
   MUX2_X1 i_132_0_436 (.A(\o_buffer[31] [11]), .B(i_mem_data[11]), .S(n_88), 
      .Z(n_132_523));
   MUX2_X1 i_132_0_437 (.A(\o_buffer[31] [10]), .B(i_mem_data[10]), .S(n_88), 
      .Z(n_132_522));
   MUX2_X1 i_132_0_438 (.A(\o_buffer[31] [9]), .B(i_mem_data[9]), .S(n_88), 
      .Z(n_132_521));
   MUX2_X1 i_132_0_439 (.A(\o_buffer[31] [8]), .B(i_mem_data[8]), .S(n_88), 
      .Z(n_132_520));
   MUX2_X1 i_132_0_440 (.A(\o_buffer[31] [7]), .B(i_mem_data[7]), .S(n_88), 
      .Z(n_132_519));
   MUX2_X1 i_132_0_441 (.A(\o_buffer[31] [6]), .B(i_mem_data[6]), .S(n_88), 
      .Z(n_132_518));
   MUX2_X1 i_132_0_442 (.A(\o_buffer[31] [5]), .B(i_mem_data[5]), .S(n_88), 
      .Z(n_132_517));
   MUX2_X1 i_132_0_443 (.A(\o_buffer[31] [4]), .B(i_mem_data[4]), .S(n_88), 
      .Z(n_132_516));
   MUX2_X1 i_132_0_444 (.A(\o_buffer[31] [3]), .B(i_mem_data[3]), .S(n_88), 
      .Z(n_132_515));
   MUX2_X1 i_132_0_445 (.A(\o_buffer[31] [2]), .B(i_mem_data[2]), .S(n_88), 
      .Z(n_132_514));
   MUX2_X1 i_132_0_446 (.A(\o_buffer[31] [1]), .B(i_mem_data[1]), .S(n_88), 
      .Z(n_132_513));
   MUX2_X1 i_132_0_447 (.A(\o_buffer[31] [0]), .B(i_mem_data[0]), .S(n_88), 
      .Z(n_132_512));
   MUX2_X1 i_132_0_448 (.A(\o_buffer[30] [15]), .B(i_mem_data[15]), .S(n_89), 
      .Z(n_132_511));
   MUX2_X1 i_132_0_449 (.A(\o_buffer[30] [14]), .B(i_mem_data[14]), .S(n_89), 
      .Z(n_132_510));
   MUX2_X1 i_132_0_450 (.A(\o_buffer[30] [13]), .B(i_mem_data[13]), .S(n_89), 
      .Z(n_132_509));
   MUX2_X1 i_132_0_451 (.A(\o_buffer[30] [12]), .B(i_mem_data[12]), .S(n_89), 
      .Z(n_132_508));
   MUX2_X1 i_132_0_452 (.A(\o_buffer[30] [11]), .B(i_mem_data[11]), .S(n_89), 
      .Z(n_132_507));
   MUX2_X1 i_132_0_453 (.A(\o_buffer[30] [10]), .B(i_mem_data[10]), .S(n_89), 
      .Z(n_132_506));
   MUX2_X1 i_132_0_454 (.A(\o_buffer[30] [9]), .B(i_mem_data[9]), .S(n_89), 
      .Z(n_132_505));
   MUX2_X1 i_132_0_455 (.A(\o_buffer[30] [8]), .B(i_mem_data[8]), .S(n_89), 
      .Z(n_132_504));
   MUX2_X1 i_132_0_456 (.A(\o_buffer[30] [7]), .B(i_mem_data[7]), .S(n_89), 
      .Z(n_132_503));
   MUX2_X1 i_132_0_457 (.A(\o_buffer[30] [6]), .B(i_mem_data[6]), .S(n_89), 
      .Z(n_132_502));
   MUX2_X1 i_132_0_458 (.A(\o_buffer[30] [5]), .B(i_mem_data[5]), .S(n_89), 
      .Z(n_132_501));
   MUX2_X1 i_132_0_459 (.A(\o_buffer[30] [4]), .B(i_mem_data[4]), .S(n_89), 
      .Z(n_132_500));
   MUX2_X1 i_132_0_460 (.A(\o_buffer[30] [3]), .B(i_mem_data[3]), .S(n_89), 
      .Z(n_132_499));
   MUX2_X1 i_132_0_461 (.A(\o_buffer[30] [2]), .B(i_mem_data[2]), .S(n_89), 
      .Z(n_132_498));
   MUX2_X1 i_132_0_462 (.A(\o_buffer[30] [1]), .B(i_mem_data[1]), .S(n_89), 
      .Z(n_132_497));
   MUX2_X1 i_132_0_463 (.A(\o_buffer[30] [0]), .B(i_mem_data[0]), .S(n_89), 
      .Z(n_132_496));
   MUX2_X1 i_132_0_464 (.A(\o_buffer[29] [15]), .B(i_mem_data[15]), .S(n_90), 
      .Z(n_132_495));
   MUX2_X1 i_132_0_465 (.A(\o_buffer[29] [14]), .B(i_mem_data[14]), .S(n_90), 
      .Z(n_132_494));
   MUX2_X1 i_132_0_466 (.A(\o_buffer[29] [13]), .B(i_mem_data[13]), .S(n_90), 
      .Z(n_132_493));
   MUX2_X1 i_132_0_467 (.A(\o_buffer[29] [12]), .B(i_mem_data[12]), .S(n_90), 
      .Z(n_132_492));
   MUX2_X1 i_132_0_468 (.A(\o_buffer[29] [11]), .B(i_mem_data[11]), .S(n_90), 
      .Z(n_132_491));
   MUX2_X1 i_132_0_469 (.A(\o_buffer[29] [10]), .B(i_mem_data[10]), .S(n_90), 
      .Z(n_132_490));
   MUX2_X1 i_132_0_470 (.A(\o_buffer[29] [9]), .B(i_mem_data[9]), .S(n_90), 
      .Z(n_132_489));
   MUX2_X1 i_132_0_471 (.A(\o_buffer[29] [8]), .B(i_mem_data[8]), .S(n_90), 
      .Z(n_132_488));
   MUX2_X1 i_132_0_472 (.A(\o_buffer[29] [7]), .B(i_mem_data[7]), .S(n_90), 
      .Z(n_132_487));
   MUX2_X1 i_132_0_473 (.A(\o_buffer[29] [6]), .B(i_mem_data[6]), .S(n_90), 
      .Z(n_132_486));
   MUX2_X1 i_132_0_474 (.A(\o_buffer[29] [5]), .B(i_mem_data[5]), .S(n_90), 
      .Z(n_132_485));
   MUX2_X1 i_132_0_475 (.A(\o_buffer[29] [4]), .B(i_mem_data[4]), .S(n_90), 
      .Z(n_132_484));
   MUX2_X1 i_132_0_476 (.A(\o_buffer[29] [3]), .B(i_mem_data[3]), .S(n_90), 
      .Z(n_132_483));
   MUX2_X1 i_132_0_477 (.A(\o_buffer[29] [2]), .B(i_mem_data[2]), .S(n_90), 
      .Z(n_132_482));
   MUX2_X1 i_132_0_478 (.A(\o_buffer[29] [1]), .B(i_mem_data[1]), .S(n_90), 
      .Z(n_132_481));
   MUX2_X1 i_132_0_479 (.A(\o_buffer[29] [0]), .B(i_mem_data[0]), .S(n_90), 
      .Z(n_132_480));
   MUX2_X1 i_132_0_480 (.A(\o_buffer[28] [15]), .B(i_mem_data[15]), .S(n_91), 
      .Z(n_132_479));
   MUX2_X1 i_132_0_481 (.A(\o_buffer[28] [14]), .B(i_mem_data[14]), .S(n_91), 
      .Z(n_132_478));
   MUX2_X1 i_132_0_482 (.A(\o_buffer[28] [13]), .B(i_mem_data[13]), .S(n_91), 
      .Z(n_132_477));
   MUX2_X1 i_132_0_483 (.A(\o_buffer[28] [12]), .B(i_mem_data[12]), .S(n_91), 
      .Z(n_132_476));
   MUX2_X1 i_132_0_484 (.A(\o_buffer[28] [11]), .B(i_mem_data[11]), .S(n_91), 
      .Z(n_132_475));
   MUX2_X1 i_132_0_485 (.A(\o_buffer[28] [10]), .B(i_mem_data[10]), .S(n_91), 
      .Z(n_132_474));
   MUX2_X1 i_132_0_486 (.A(\o_buffer[28] [9]), .B(i_mem_data[9]), .S(n_91), 
      .Z(n_132_473));
   MUX2_X1 i_132_0_487 (.A(\o_buffer[28] [8]), .B(i_mem_data[8]), .S(n_91), 
      .Z(n_132_472));
   MUX2_X1 i_132_0_488 (.A(\o_buffer[28] [7]), .B(i_mem_data[7]), .S(n_91), 
      .Z(n_132_471));
   MUX2_X1 i_132_0_489 (.A(\o_buffer[28] [6]), .B(i_mem_data[6]), .S(n_91), 
      .Z(n_132_470));
   MUX2_X1 i_132_0_490 (.A(\o_buffer[28] [5]), .B(i_mem_data[5]), .S(n_91), 
      .Z(n_132_469));
   MUX2_X1 i_132_0_491 (.A(\o_buffer[28] [4]), .B(i_mem_data[4]), .S(n_91), 
      .Z(n_132_468));
   MUX2_X1 i_132_0_492 (.A(\o_buffer[28] [3]), .B(i_mem_data[3]), .S(n_91), 
      .Z(n_132_467));
   MUX2_X1 i_132_0_493 (.A(\o_buffer[28] [2]), .B(i_mem_data[2]), .S(n_91), 
      .Z(n_132_466));
   MUX2_X1 i_132_0_494 (.A(\o_buffer[28] [1]), .B(i_mem_data[1]), .S(n_91), 
      .Z(n_132_465));
   MUX2_X1 i_132_0_495 (.A(\o_buffer[28] [0]), .B(i_mem_data[0]), .S(n_91), 
      .Z(n_132_464));
   MUX2_X1 i_132_0_496 (.A(\o_buffer[27] [15]), .B(i_mem_data[15]), .S(n_92), 
      .Z(n_132_463));
   MUX2_X1 i_132_0_497 (.A(\o_buffer[27] [14]), .B(i_mem_data[14]), .S(n_92), 
      .Z(n_132_462));
   MUX2_X1 i_132_0_498 (.A(\o_buffer[27] [13]), .B(i_mem_data[13]), .S(n_92), 
      .Z(n_132_461));
   MUX2_X1 i_132_0_499 (.A(\o_buffer[27] [12]), .B(i_mem_data[12]), .S(n_92), 
      .Z(n_132_460));
   MUX2_X1 i_132_0_500 (.A(\o_buffer[27] [11]), .B(i_mem_data[11]), .S(n_92), 
      .Z(n_132_459));
   MUX2_X1 i_132_0_501 (.A(\o_buffer[27] [10]), .B(i_mem_data[10]), .S(n_92), 
      .Z(n_132_458));
   MUX2_X1 i_132_0_502 (.A(\o_buffer[27] [9]), .B(i_mem_data[9]), .S(n_92), 
      .Z(n_132_457));
   MUX2_X1 i_132_0_503 (.A(\o_buffer[27] [8]), .B(i_mem_data[8]), .S(n_92), 
      .Z(n_132_456));
   MUX2_X1 i_132_0_504 (.A(\o_buffer[27] [7]), .B(i_mem_data[7]), .S(n_92), 
      .Z(n_132_455));
   MUX2_X1 i_132_0_505 (.A(\o_buffer[27] [6]), .B(i_mem_data[6]), .S(n_92), 
      .Z(n_132_454));
   MUX2_X1 i_132_0_506 (.A(\o_buffer[27] [5]), .B(i_mem_data[5]), .S(n_92), 
      .Z(n_132_453));
   MUX2_X1 i_132_0_507 (.A(\o_buffer[27] [4]), .B(i_mem_data[4]), .S(n_92), 
      .Z(n_132_452));
   MUX2_X1 i_132_0_508 (.A(\o_buffer[27] [3]), .B(i_mem_data[3]), .S(n_92), 
      .Z(n_132_451));
   MUX2_X1 i_132_0_509 (.A(\o_buffer[27] [2]), .B(i_mem_data[2]), .S(n_92), 
      .Z(n_132_450));
   MUX2_X1 i_132_0_510 (.A(\o_buffer[27] [1]), .B(i_mem_data[1]), .S(n_92), 
      .Z(n_132_449));
   MUX2_X1 i_132_0_511 (.A(\o_buffer[27] [0]), .B(i_mem_data[0]), .S(n_92), 
      .Z(n_132_448));
   MUX2_X1 i_132_0_512 (.A(\o_buffer[26] [15]), .B(i_mem_data[15]), .S(n_93), 
      .Z(n_132_447));
   MUX2_X1 i_132_0_513 (.A(\o_buffer[26] [14]), .B(i_mem_data[14]), .S(n_93), 
      .Z(n_132_446));
   MUX2_X1 i_132_0_514 (.A(\o_buffer[26] [13]), .B(i_mem_data[13]), .S(n_93), 
      .Z(n_132_445));
   MUX2_X1 i_132_0_515 (.A(\o_buffer[26] [12]), .B(i_mem_data[12]), .S(n_93), 
      .Z(n_132_444));
   MUX2_X1 i_132_0_516 (.A(\o_buffer[26] [11]), .B(i_mem_data[11]), .S(n_93), 
      .Z(n_132_443));
   MUX2_X1 i_132_0_517 (.A(\o_buffer[26] [10]), .B(i_mem_data[10]), .S(n_93), 
      .Z(n_132_442));
   MUX2_X1 i_132_0_518 (.A(\o_buffer[26] [9]), .B(i_mem_data[9]), .S(n_93), 
      .Z(n_132_441));
   MUX2_X1 i_132_0_519 (.A(\o_buffer[26] [8]), .B(i_mem_data[8]), .S(n_93), 
      .Z(n_132_440));
   MUX2_X1 i_132_0_520 (.A(\o_buffer[26] [7]), .B(i_mem_data[7]), .S(n_93), 
      .Z(n_132_439));
   MUX2_X1 i_132_0_521 (.A(\o_buffer[26] [6]), .B(i_mem_data[6]), .S(n_93), 
      .Z(n_132_438));
   MUX2_X1 i_132_0_522 (.A(\o_buffer[26] [5]), .B(i_mem_data[5]), .S(n_93), 
      .Z(n_132_437));
   MUX2_X1 i_132_0_523 (.A(\o_buffer[26] [4]), .B(i_mem_data[4]), .S(n_93), 
      .Z(n_132_436));
   MUX2_X1 i_132_0_524 (.A(\o_buffer[26] [3]), .B(i_mem_data[3]), .S(n_93), 
      .Z(n_132_435));
   MUX2_X1 i_132_0_525 (.A(\o_buffer[26] [2]), .B(i_mem_data[2]), .S(n_93), 
      .Z(n_132_434));
   MUX2_X1 i_132_0_526 (.A(\o_buffer[26] [1]), .B(i_mem_data[1]), .S(n_93), 
      .Z(n_132_433));
   MUX2_X1 i_132_0_527 (.A(\o_buffer[26] [0]), .B(i_mem_data[0]), .S(n_93), 
      .Z(n_132_432));
   MUX2_X1 i_132_0_528 (.A(\o_buffer[25] [15]), .B(i_mem_data[15]), .S(n_94), 
      .Z(n_132_431));
   MUX2_X1 i_132_0_529 (.A(\o_buffer[25] [14]), .B(i_mem_data[14]), .S(n_94), 
      .Z(n_132_430));
   MUX2_X1 i_132_0_530 (.A(\o_buffer[25] [13]), .B(i_mem_data[13]), .S(n_94), 
      .Z(n_132_429));
   MUX2_X1 i_132_0_531 (.A(\o_buffer[25] [12]), .B(i_mem_data[12]), .S(n_94), 
      .Z(n_132_428));
   MUX2_X1 i_132_0_532 (.A(\o_buffer[25] [11]), .B(i_mem_data[11]), .S(n_94), 
      .Z(n_132_427));
   MUX2_X1 i_132_0_533 (.A(\o_buffer[25] [10]), .B(i_mem_data[10]), .S(n_94), 
      .Z(n_132_426));
   MUX2_X1 i_132_0_534 (.A(\o_buffer[25] [9]), .B(i_mem_data[9]), .S(n_94), 
      .Z(n_132_425));
   MUX2_X1 i_132_0_535 (.A(\o_buffer[25] [8]), .B(i_mem_data[8]), .S(n_94), 
      .Z(n_132_424));
   MUX2_X1 i_132_0_536 (.A(\o_buffer[25] [7]), .B(i_mem_data[7]), .S(n_94), 
      .Z(n_132_423));
   MUX2_X1 i_132_0_537 (.A(\o_buffer[25] [6]), .B(i_mem_data[6]), .S(n_94), 
      .Z(n_132_422));
   MUX2_X1 i_132_0_538 (.A(\o_buffer[25] [5]), .B(i_mem_data[5]), .S(n_94), 
      .Z(n_132_421));
   MUX2_X1 i_132_0_539 (.A(\o_buffer[25] [4]), .B(i_mem_data[4]), .S(n_94), 
      .Z(n_132_420));
   MUX2_X1 i_132_0_540 (.A(\o_buffer[25] [3]), .B(i_mem_data[3]), .S(n_94), 
      .Z(n_132_419));
   MUX2_X1 i_132_0_541 (.A(\o_buffer[25] [2]), .B(i_mem_data[2]), .S(n_94), 
      .Z(n_132_418));
   MUX2_X1 i_132_0_542 (.A(\o_buffer[25] [1]), .B(i_mem_data[1]), .S(n_94), 
      .Z(n_132_417));
   MUX2_X1 i_132_0_543 (.A(\o_buffer[25] [0]), .B(i_mem_data[0]), .S(n_94), 
      .Z(n_132_416));
   MUX2_X1 i_132_0_544 (.A(\o_buffer[24] [15]), .B(i_mem_data[15]), .S(n_95), 
      .Z(n_132_415));
   MUX2_X1 i_132_0_545 (.A(\o_buffer[24] [14]), .B(i_mem_data[14]), .S(n_95), 
      .Z(n_132_414));
   MUX2_X1 i_132_0_546 (.A(\o_buffer[24] [13]), .B(i_mem_data[13]), .S(n_95), 
      .Z(n_132_413));
   MUX2_X1 i_132_0_547 (.A(\o_buffer[24] [12]), .B(i_mem_data[12]), .S(n_95), 
      .Z(n_132_412));
   MUX2_X1 i_132_0_548 (.A(\o_buffer[24] [11]), .B(i_mem_data[11]), .S(n_95), 
      .Z(n_132_411));
   MUX2_X1 i_132_0_549 (.A(\o_buffer[24] [10]), .B(i_mem_data[10]), .S(n_95), 
      .Z(n_132_410));
   MUX2_X1 i_132_0_550 (.A(\o_buffer[24] [9]), .B(i_mem_data[9]), .S(n_95), 
      .Z(n_132_409));
   MUX2_X1 i_132_0_551 (.A(\o_buffer[24] [8]), .B(i_mem_data[8]), .S(n_95), 
      .Z(n_132_408));
   MUX2_X1 i_132_0_552 (.A(\o_buffer[24] [7]), .B(i_mem_data[7]), .S(n_95), 
      .Z(n_132_407));
   MUX2_X1 i_132_0_553 (.A(\o_buffer[24] [6]), .B(i_mem_data[6]), .S(n_95), 
      .Z(n_132_406));
   MUX2_X1 i_132_0_554 (.A(\o_buffer[24] [5]), .B(i_mem_data[5]), .S(n_95), 
      .Z(n_132_405));
   MUX2_X1 i_132_0_555 (.A(\o_buffer[24] [4]), .B(i_mem_data[4]), .S(n_95), 
      .Z(n_132_404));
   MUX2_X1 i_132_0_556 (.A(\o_buffer[24] [3]), .B(i_mem_data[3]), .S(n_95), 
      .Z(n_132_403));
   MUX2_X1 i_132_0_557 (.A(\o_buffer[24] [2]), .B(i_mem_data[2]), .S(n_95), 
      .Z(n_132_402));
   MUX2_X1 i_132_0_558 (.A(\o_buffer[24] [1]), .B(i_mem_data[1]), .S(n_95), 
      .Z(n_132_401));
   MUX2_X1 i_132_0_559 (.A(\o_buffer[24] [0]), .B(i_mem_data[0]), .S(n_95), 
      .Z(n_132_400));
   MUX2_X1 i_132_0_560 (.A(\o_buffer[23] [15]), .B(i_mem_data[15]), .S(n_96), 
      .Z(n_132_399));
   MUX2_X1 i_132_0_561 (.A(\o_buffer[23] [14]), .B(i_mem_data[14]), .S(n_96), 
      .Z(n_132_398));
   MUX2_X1 i_132_0_562 (.A(\o_buffer[23] [13]), .B(i_mem_data[13]), .S(n_96), 
      .Z(n_132_397));
   MUX2_X1 i_132_0_563 (.A(\o_buffer[23] [12]), .B(i_mem_data[12]), .S(n_96), 
      .Z(n_132_396));
   MUX2_X1 i_132_0_564 (.A(\o_buffer[23] [11]), .B(i_mem_data[11]), .S(n_96), 
      .Z(n_132_395));
   MUX2_X1 i_132_0_565 (.A(\o_buffer[23] [10]), .B(i_mem_data[10]), .S(n_96), 
      .Z(n_132_394));
   MUX2_X1 i_132_0_566 (.A(\o_buffer[23] [9]), .B(i_mem_data[9]), .S(n_96), 
      .Z(n_132_393));
   MUX2_X1 i_132_0_567 (.A(\o_buffer[23] [8]), .B(i_mem_data[8]), .S(n_96), 
      .Z(n_132_392));
   MUX2_X1 i_132_0_568 (.A(\o_buffer[23] [7]), .B(i_mem_data[7]), .S(n_96), 
      .Z(n_132_391));
   MUX2_X1 i_132_0_569 (.A(\o_buffer[23] [6]), .B(i_mem_data[6]), .S(n_96), 
      .Z(n_132_390));
   MUX2_X1 i_132_0_570 (.A(\o_buffer[23] [5]), .B(i_mem_data[5]), .S(n_96), 
      .Z(n_132_389));
   MUX2_X1 i_132_0_571 (.A(\o_buffer[23] [4]), .B(i_mem_data[4]), .S(n_96), 
      .Z(n_132_388));
   MUX2_X1 i_132_0_572 (.A(\o_buffer[23] [3]), .B(i_mem_data[3]), .S(n_96), 
      .Z(n_132_387));
   MUX2_X1 i_132_0_573 (.A(\o_buffer[23] [2]), .B(i_mem_data[2]), .S(n_96), 
      .Z(n_132_386));
   MUX2_X1 i_132_0_574 (.A(\o_buffer[23] [1]), .B(i_mem_data[1]), .S(n_96), 
      .Z(n_132_385));
   MUX2_X1 i_132_0_575 (.A(\o_buffer[23] [0]), .B(i_mem_data[0]), .S(n_96), 
      .Z(n_132_384));
   MUX2_X1 i_132_0_576 (.A(\o_buffer[22] [15]), .B(i_mem_data[15]), .S(n_97), 
      .Z(n_132_383));
   MUX2_X1 i_132_0_577 (.A(\o_buffer[22] [14]), .B(i_mem_data[14]), .S(n_97), 
      .Z(n_132_382));
   MUX2_X1 i_132_0_578 (.A(\o_buffer[22] [13]), .B(i_mem_data[13]), .S(n_97), 
      .Z(n_132_381));
   MUX2_X1 i_132_0_579 (.A(\o_buffer[22] [12]), .B(i_mem_data[12]), .S(n_97), 
      .Z(n_132_380));
   MUX2_X1 i_132_0_580 (.A(\o_buffer[22] [11]), .B(i_mem_data[11]), .S(n_97), 
      .Z(n_132_379));
   MUX2_X1 i_132_0_581 (.A(\o_buffer[22] [10]), .B(i_mem_data[10]), .S(n_97), 
      .Z(n_132_378));
   MUX2_X1 i_132_0_582 (.A(\o_buffer[22] [9]), .B(i_mem_data[9]), .S(n_97), 
      .Z(n_132_377));
   MUX2_X1 i_132_0_583 (.A(\o_buffer[22] [8]), .B(i_mem_data[8]), .S(n_97), 
      .Z(n_132_376));
   MUX2_X1 i_132_0_584 (.A(\o_buffer[22] [7]), .B(i_mem_data[7]), .S(n_97), 
      .Z(n_132_375));
   MUX2_X1 i_132_0_585 (.A(\o_buffer[22] [6]), .B(i_mem_data[6]), .S(n_97), 
      .Z(n_132_374));
   MUX2_X1 i_132_0_586 (.A(\o_buffer[22] [5]), .B(i_mem_data[5]), .S(n_97), 
      .Z(n_132_373));
   MUX2_X1 i_132_0_587 (.A(\o_buffer[22] [4]), .B(i_mem_data[4]), .S(n_97), 
      .Z(n_132_372));
   MUX2_X1 i_132_0_588 (.A(\o_buffer[22] [3]), .B(i_mem_data[3]), .S(n_97), 
      .Z(n_132_371));
   MUX2_X1 i_132_0_589 (.A(\o_buffer[22] [2]), .B(i_mem_data[2]), .S(n_97), 
      .Z(n_132_370));
   MUX2_X1 i_132_0_590 (.A(\o_buffer[22] [1]), .B(i_mem_data[1]), .S(n_97), 
      .Z(n_132_369));
   MUX2_X1 i_132_0_591 (.A(\o_buffer[22] [0]), .B(i_mem_data[0]), .S(n_97), 
      .Z(n_132_368));
   MUX2_X1 i_132_0_592 (.A(\o_buffer[21] [15]), .B(i_mem_data[15]), .S(n_98), 
      .Z(n_132_367));
   MUX2_X1 i_132_0_593 (.A(\o_buffer[21] [14]), .B(i_mem_data[14]), .S(n_98), 
      .Z(n_132_366));
   MUX2_X1 i_132_0_594 (.A(\o_buffer[21] [13]), .B(i_mem_data[13]), .S(n_98), 
      .Z(n_132_365));
   MUX2_X1 i_132_0_595 (.A(\o_buffer[21] [12]), .B(i_mem_data[12]), .S(n_98), 
      .Z(n_132_364));
   MUX2_X1 i_132_0_596 (.A(\o_buffer[21] [11]), .B(i_mem_data[11]), .S(n_98), 
      .Z(n_132_363));
   MUX2_X1 i_132_0_597 (.A(\o_buffer[21] [10]), .B(i_mem_data[10]), .S(n_98), 
      .Z(n_132_362));
   MUX2_X1 i_132_0_598 (.A(\o_buffer[21] [9]), .B(i_mem_data[9]), .S(n_98), 
      .Z(n_132_361));
   MUX2_X1 i_132_0_599 (.A(\o_buffer[21] [8]), .B(i_mem_data[8]), .S(n_98), 
      .Z(n_132_360));
   MUX2_X1 i_132_0_600 (.A(\o_buffer[21] [7]), .B(i_mem_data[7]), .S(n_98), 
      .Z(n_132_359));
   MUX2_X1 i_132_0_601 (.A(\o_buffer[21] [6]), .B(i_mem_data[6]), .S(n_98), 
      .Z(n_132_358));
   MUX2_X1 i_132_0_602 (.A(\o_buffer[21] [5]), .B(i_mem_data[5]), .S(n_98), 
      .Z(n_132_357));
   MUX2_X1 i_132_0_603 (.A(\o_buffer[21] [4]), .B(i_mem_data[4]), .S(n_98), 
      .Z(n_132_356));
   MUX2_X1 i_132_0_604 (.A(\o_buffer[21] [3]), .B(i_mem_data[3]), .S(n_98), 
      .Z(n_132_355));
   MUX2_X1 i_132_0_605 (.A(\o_buffer[21] [2]), .B(i_mem_data[2]), .S(n_98), 
      .Z(n_132_354));
   MUX2_X1 i_132_0_606 (.A(\o_buffer[21] [1]), .B(i_mem_data[1]), .S(n_98), 
      .Z(n_132_353));
   MUX2_X1 i_132_0_607 (.A(\o_buffer[21] [0]), .B(i_mem_data[0]), .S(n_98), 
      .Z(n_132_352));
   MUX2_X1 i_132_0_608 (.A(\o_buffer[20] [15]), .B(i_mem_data[15]), .S(n_99), 
      .Z(n_132_351));
   MUX2_X1 i_132_0_609 (.A(\o_buffer[20] [14]), .B(i_mem_data[14]), .S(n_99), 
      .Z(n_132_350));
   MUX2_X1 i_132_0_610 (.A(\o_buffer[20] [13]), .B(i_mem_data[13]), .S(n_99), 
      .Z(n_132_349));
   MUX2_X1 i_132_0_611 (.A(\o_buffer[20] [12]), .B(i_mem_data[12]), .S(n_99), 
      .Z(n_132_348));
   MUX2_X1 i_132_0_612 (.A(\o_buffer[20] [11]), .B(i_mem_data[11]), .S(n_99), 
      .Z(n_132_347));
   MUX2_X1 i_132_0_613 (.A(\o_buffer[20] [10]), .B(i_mem_data[10]), .S(n_99), 
      .Z(n_132_346));
   MUX2_X1 i_132_0_614 (.A(\o_buffer[20] [9]), .B(i_mem_data[9]), .S(n_99), 
      .Z(n_132_345));
   MUX2_X1 i_132_0_615 (.A(\o_buffer[20] [8]), .B(i_mem_data[8]), .S(n_99), 
      .Z(n_132_344));
   MUX2_X1 i_132_0_616 (.A(\o_buffer[20] [7]), .B(i_mem_data[7]), .S(n_99), 
      .Z(n_132_343));
   MUX2_X1 i_132_0_617 (.A(\o_buffer[20] [6]), .B(i_mem_data[6]), .S(n_99), 
      .Z(n_132_342));
   MUX2_X1 i_132_0_618 (.A(\o_buffer[20] [5]), .B(i_mem_data[5]), .S(n_99), 
      .Z(n_132_341));
   MUX2_X1 i_132_0_619 (.A(\o_buffer[20] [4]), .B(i_mem_data[4]), .S(n_99), 
      .Z(n_132_340));
   MUX2_X1 i_132_0_620 (.A(\o_buffer[20] [3]), .B(i_mem_data[3]), .S(n_99), 
      .Z(n_132_339));
   MUX2_X1 i_132_0_621 (.A(\o_buffer[20] [2]), .B(i_mem_data[2]), .S(n_99), 
      .Z(n_132_338));
   MUX2_X1 i_132_0_622 (.A(\o_buffer[20] [1]), .B(i_mem_data[1]), .S(n_99), 
      .Z(n_132_337));
   MUX2_X1 i_132_0_623 (.A(\o_buffer[20] [0]), .B(i_mem_data[0]), .S(n_99), 
      .Z(n_132_336));
   MUX2_X1 i_132_0_624 (.A(\o_buffer[19] [15]), .B(i_mem_data[15]), .S(n_100), 
      .Z(n_132_335));
   MUX2_X1 i_132_0_625 (.A(\o_buffer[19] [14]), .B(i_mem_data[14]), .S(n_100), 
      .Z(n_132_334));
   MUX2_X1 i_132_0_626 (.A(\o_buffer[19] [13]), .B(i_mem_data[13]), .S(n_100), 
      .Z(n_132_333));
   MUX2_X1 i_132_0_627 (.A(\o_buffer[19] [12]), .B(i_mem_data[12]), .S(n_100), 
      .Z(n_132_332));
   MUX2_X1 i_132_0_628 (.A(\o_buffer[19] [11]), .B(i_mem_data[11]), .S(n_100), 
      .Z(n_132_331));
   MUX2_X1 i_132_0_629 (.A(\o_buffer[19] [10]), .B(i_mem_data[10]), .S(n_100), 
      .Z(n_132_330));
   MUX2_X1 i_132_0_630 (.A(\o_buffer[19] [9]), .B(i_mem_data[9]), .S(n_100), 
      .Z(n_132_329));
   MUX2_X1 i_132_0_631 (.A(\o_buffer[19] [8]), .B(i_mem_data[8]), .S(n_100), 
      .Z(n_132_328));
   MUX2_X1 i_132_0_632 (.A(\o_buffer[19] [7]), .B(i_mem_data[7]), .S(n_100), 
      .Z(n_132_327));
   MUX2_X1 i_132_0_633 (.A(\o_buffer[19] [6]), .B(i_mem_data[6]), .S(n_100), 
      .Z(n_132_326));
   MUX2_X1 i_132_0_634 (.A(\o_buffer[19] [5]), .B(i_mem_data[5]), .S(n_100), 
      .Z(n_132_325));
   MUX2_X1 i_132_0_635 (.A(\o_buffer[19] [4]), .B(i_mem_data[4]), .S(n_100), 
      .Z(n_132_324));
   MUX2_X1 i_132_0_636 (.A(\o_buffer[19] [3]), .B(i_mem_data[3]), .S(n_100), 
      .Z(n_132_323));
   MUX2_X1 i_132_0_637 (.A(\o_buffer[19] [2]), .B(i_mem_data[2]), .S(n_100), 
      .Z(n_132_322));
   MUX2_X1 i_132_0_638 (.A(\o_buffer[19] [1]), .B(i_mem_data[1]), .S(n_100), 
      .Z(n_132_321));
   MUX2_X1 i_132_0_639 (.A(\o_buffer[19] [0]), .B(i_mem_data[0]), .S(n_100), 
      .Z(n_132_320));
   MUX2_X1 i_132_0_640 (.A(\o_buffer[18] [15]), .B(i_mem_data[15]), .S(n_101), 
      .Z(n_132_319));
   MUX2_X1 i_132_0_641 (.A(\o_buffer[18] [14]), .B(i_mem_data[14]), .S(n_101), 
      .Z(n_132_318));
   MUX2_X1 i_132_0_642 (.A(\o_buffer[18] [13]), .B(i_mem_data[13]), .S(n_101), 
      .Z(n_132_317));
   MUX2_X1 i_132_0_643 (.A(\o_buffer[18] [12]), .B(i_mem_data[12]), .S(n_101), 
      .Z(n_132_316));
   MUX2_X1 i_132_0_644 (.A(\o_buffer[18] [11]), .B(i_mem_data[11]), .S(n_101), 
      .Z(n_132_315));
   MUX2_X1 i_132_0_645 (.A(\o_buffer[18] [10]), .B(i_mem_data[10]), .S(n_101), 
      .Z(n_132_314));
   MUX2_X1 i_132_0_646 (.A(\o_buffer[18] [9]), .B(i_mem_data[9]), .S(n_101), 
      .Z(n_132_313));
   MUX2_X1 i_132_0_647 (.A(\o_buffer[18] [8]), .B(i_mem_data[8]), .S(n_101), 
      .Z(n_132_312));
   MUX2_X1 i_132_0_648 (.A(\o_buffer[18] [7]), .B(i_mem_data[7]), .S(n_101), 
      .Z(n_132_311));
   MUX2_X1 i_132_0_649 (.A(\o_buffer[18] [6]), .B(i_mem_data[6]), .S(n_101), 
      .Z(n_132_310));
   MUX2_X1 i_132_0_650 (.A(\o_buffer[18] [5]), .B(i_mem_data[5]), .S(n_101), 
      .Z(n_132_309));
   MUX2_X1 i_132_0_651 (.A(\o_buffer[18] [4]), .B(i_mem_data[4]), .S(n_101), 
      .Z(n_132_308));
   MUX2_X1 i_132_0_652 (.A(\o_buffer[18] [3]), .B(i_mem_data[3]), .S(n_101), 
      .Z(n_132_307));
   MUX2_X1 i_132_0_653 (.A(\o_buffer[18] [2]), .B(i_mem_data[2]), .S(n_101), 
      .Z(n_132_306));
   MUX2_X1 i_132_0_654 (.A(\o_buffer[18] [1]), .B(i_mem_data[1]), .S(n_101), 
      .Z(n_132_305));
   MUX2_X1 i_132_0_655 (.A(\o_buffer[18] [0]), .B(i_mem_data[0]), .S(n_101), 
      .Z(n_132_304));
   MUX2_X1 i_132_0_656 (.A(\o_buffer[17] [15]), .B(i_mem_data[15]), .S(n_102), 
      .Z(n_132_303));
   MUX2_X1 i_132_0_657 (.A(\o_buffer[17] [14]), .B(i_mem_data[14]), .S(n_102), 
      .Z(n_132_302));
   MUX2_X1 i_132_0_658 (.A(\o_buffer[17] [13]), .B(i_mem_data[13]), .S(n_102), 
      .Z(n_132_301));
   MUX2_X1 i_132_0_659 (.A(\o_buffer[17] [12]), .B(i_mem_data[12]), .S(n_102), 
      .Z(n_132_300));
   MUX2_X1 i_132_0_660 (.A(\o_buffer[17] [11]), .B(i_mem_data[11]), .S(n_102), 
      .Z(n_132_299));
   MUX2_X1 i_132_0_661 (.A(\o_buffer[17] [10]), .B(i_mem_data[10]), .S(n_102), 
      .Z(n_132_298));
   MUX2_X1 i_132_0_662 (.A(\o_buffer[17] [9]), .B(i_mem_data[9]), .S(n_102), 
      .Z(n_132_297));
   MUX2_X1 i_132_0_663 (.A(\o_buffer[17] [8]), .B(i_mem_data[8]), .S(n_102), 
      .Z(n_132_296));
   MUX2_X1 i_132_0_664 (.A(\o_buffer[17] [7]), .B(i_mem_data[7]), .S(n_102), 
      .Z(n_132_295));
   MUX2_X1 i_132_0_665 (.A(\o_buffer[17] [6]), .B(i_mem_data[6]), .S(n_102), 
      .Z(n_132_294));
   MUX2_X1 i_132_0_666 (.A(\o_buffer[17] [5]), .B(i_mem_data[5]), .S(n_102), 
      .Z(n_132_293));
   MUX2_X1 i_132_0_667 (.A(\o_buffer[17] [4]), .B(i_mem_data[4]), .S(n_102), 
      .Z(n_132_292));
   MUX2_X1 i_132_0_668 (.A(\o_buffer[17] [3]), .B(i_mem_data[3]), .S(n_102), 
      .Z(n_132_291));
   MUX2_X1 i_132_0_669 (.A(\o_buffer[17] [2]), .B(i_mem_data[2]), .S(n_102), 
      .Z(n_132_290));
   MUX2_X1 i_132_0_670 (.A(\o_buffer[17] [1]), .B(i_mem_data[1]), .S(n_102), 
      .Z(n_132_289));
   MUX2_X1 i_132_0_671 (.A(\o_buffer[17] [0]), .B(i_mem_data[0]), .S(n_102), 
      .Z(n_132_288));
   MUX2_X1 i_132_0_672 (.A(\o_buffer[16] [15]), .B(i_mem_data[15]), .S(n_103), 
      .Z(n_132_287));
   MUX2_X1 i_132_0_673 (.A(\o_buffer[16] [14]), .B(i_mem_data[14]), .S(n_103), 
      .Z(n_132_286));
   MUX2_X1 i_132_0_674 (.A(\o_buffer[16] [13]), .B(i_mem_data[13]), .S(n_103), 
      .Z(n_132_285));
   MUX2_X1 i_132_0_675 (.A(\o_buffer[16] [12]), .B(i_mem_data[12]), .S(n_103), 
      .Z(n_132_284));
   MUX2_X1 i_132_0_676 (.A(\o_buffer[16] [11]), .B(i_mem_data[11]), .S(n_103), 
      .Z(n_132_283));
   MUX2_X1 i_132_0_677 (.A(\o_buffer[16] [10]), .B(i_mem_data[10]), .S(n_103), 
      .Z(n_132_282));
   MUX2_X1 i_132_0_678 (.A(\o_buffer[16] [9]), .B(i_mem_data[9]), .S(n_103), 
      .Z(n_132_281));
   MUX2_X1 i_132_0_679 (.A(\o_buffer[16] [8]), .B(i_mem_data[8]), .S(n_103), 
      .Z(n_132_280));
   MUX2_X1 i_132_0_680 (.A(\o_buffer[16] [7]), .B(i_mem_data[7]), .S(n_103), 
      .Z(n_132_279));
   MUX2_X1 i_132_0_681 (.A(\o_buffer[16] [6]), .B(i_mem_data[6]), .S(n_103), 
      .Z(n_132_278));
   MUX2_X1 i_132_0_682 (.A(\o_buffer[16] [5]), .B(i_mem_data[5]), .S(n_103), 
      .Z(n_132_277));
   MUX2_X1 i_132_0_683 (.A(\o_buffer[16] [4]), .B(i_mem_data[4]), .S(n_103), 
      .Z(n_132_276));
   MUX2_X1 i_132_0_684 (.A(\o_buffer[16] [3]), .B(i_mem_data[3]), .S(n_103), 
      .Z(n_132_275));
   MUX2_X1 i_132_0_685 (.A(\o_buffer[16] [2]), .B(i_mem_data[2]), .S(n_103), 
      .Z(n_132_274));
   MUX2_X1 i_132_0_686 (.A(\o_buffer[16] [1]), .B(i_mem_data[1]), .S(n_103), 
      .Z(n_132_273));
   MUX2_X1 i_132_0_687 (.A(\o_buffer[16] [0]), .B(i_mem_data[0]), .S(n_103), 
      .Z(n_132_272));
   MUX2_X1 i_132_0_688 (.A(\o_buffer[15] [15]), .B(i_mem_data[15]), .S(n_104), 
      .Z(n_132_271));
   MUX2_X1 i_132_0_689 (.A(\o_buffer[15] [14]), .B(i_mem_data[14]), .S(n_104), 
      .Z(n_132_270));
   MUX2_X1 i_132_0_690 (.A(\o_buffer[15] [13]), .B(i_mem_data[13]), .S(n_104), 
      .Z(n_132_269));
   MUX2_X1 i_132_0_691 (.A(\o_buffer[15] [12]), .B(i_mem_data[12]), .S(n_104), 
      .Z(n_132_268));
   MUX2_X1 i_132_0_692 (.A(\o_buffer[15] [11]), .B(i_mem_data[11]), .S(n_104), 
      .Z(n_132_267));
   MUX2_X1 i_132_0_693 (.A(\o_buffer[15] [10]), .B(i_mem_data[10]), .S(n_104), 
      .Z(n_132_266));
   MUX2_X1 i_132_0_694 (.A(\o_buffer[15] [9]), .B(i_mem_data[9]), .S(n_104), 
      .Z(n_132_265));
   MUX2_X1 i_132_0_695 (.A(\o_buffer[15] [8]), .B(i_mem_data[8]), .S(n_104), 
      .Z(n_132_264));
   MUX2_X1 i_132_0_696 (.A(\o_buffer[15] [7]), .B(i_mem_data[7]), .S(n_104), 
      .Z(n_132_263));
   MUX2_X1 i_132_0_697 (.A(\o_buffer[15] [6]), .B(i_mem_data[6]), .S(n_104), 
      .Z(n_132_262));
   MUX2_X1 i_132_0_698 (.A(\o_buffer[15] [5]), .B(i_mem_data[5]), .S(n_104), 
      .Z(n_132_261));
   MUX2_X1 i_132_0_699 (.A(\o_buffer[15] [4]), .B(i_mem_data[4]), .S(n_104), 
      .Z(n_132_260));
   MUX2_X1 i_132_0_700 (.A(\o_buffer[15] [3]), .B(i_mem_data[3]), .S(n_104), 
      .Z(n_132_259));
   MUX2_X1 i_132_0_701 (.A(\o_buffer[15] [2]), .B(i_mem_data[2]), .S(n_104), 
      .Z(n_132_258));
   MUX2_X1 i_132_0_702 (.A(\o_buffer[15] [1]), .B(i_mem_data[1]), .S(n_104), 
      .Z(n_132_257));
   MUX2_X1 i_132_0_703 (.A(\o_buffer[15] [0]), .B(i_mem_data[0]), .S(n_104), 
      .Z(n_132_256));
   MUX2_X1 i_132_0_704 (.A(\o_buffer[14] [15]), .B(i_mem_data[15]), .S(n_105), 
      .Z(n_132_255));
   MUX2_X1 i_132_0_705 (.A(\o_buffer[14] [14]), .B(i_mem_data[14]), .S(n_105), 
      .Z(n_132_254));
   MUX2_X1 i_132_0_706 (.A(\o_buffer[14] [13]), .B(i_mem_data[13]), .S(n_105), 
      .Z(n_132_253));
   MUX2_X1 i_132_0_707 (.A(\o_buffer[14] [12]), .B(i_mem_data[12]), .S(n_105), 
      .Z(n_132_252));
   MUX2_X1 i_132_0_708 (.A(\o_buffer[14] [11]), .B(i_mem_data[11]), .S(n_105), 
      .Z(n_132_251));
   MUX2_X1 i_132_0_709 (.A(\o_buffer[14] [10]), .B(i_mem_data[10]), .S(n_105), 
      .Z(n_132_250));
   MUX2_X1 i_132_0_710 (.A(\o_buffer[14] [9]), .B(i_mem_data[9]), .S(n_105), 
      .Z(n_132_249));
   MUX2_X1 i_132_0_711 (.A(\o_buffer[14] [8]), .B(i_mem_data[8]), .S(n_105), 
      .Z(n_132_248));
   MUX2_X1 i_132_0_712 (.A(\o_buffer[14] [7]), .B(i_mem_data[7]), .S(n_105), 
      .Z(n_132_247));
   MUX2_X1 i_132_0_713 (.A(\o_buffer[14] [6]), .B(i_mem_data[6]), .S(n_105), 
      .Z(n_132_246));
   MUX2_X1 i_132_0_714 (.A(\o_buffer[14] [5]), .B(i_mem_data[5]), .S(n_105), 
      .Z(n_132_245));
   MUX2_X1 i_132_0_715 (.A(\o_buffer[14] [4]), .B(i_mem_data[4]), .S(n_105), 
      .Z(n_132_244));
   MUX2_X1 i_132_0_716 (.A(\o_buffer[14] [3]), .B(i_mem_data[3]), .S(n_105), 
      .Z(n_132_243));
   MUX2_X1 i_132_0_717 (.A(\o_buffer[14] [2]), .B(i_mem_data[2]), .S(n_105), 
      .Z(n_132_242));
   MUX2_X1 i_132_0_718 (.A(\o_buffer[14] [1]), .B(i_mem_data[1]), .S(n_105), 
      .Z(n_132_241));
   MUX2_X1 i_132_0_719 (.A(\o_buffer[14] [0]), .B(i_mem_data[0]), .S(n_105), 
      .Z(n_132_240));
   MUX2_X1 i_132_0_720 (.A(\o_buffer[13] [15]), .B(i_mem_data[15]), .S(n_106), 
      .Z(n_132_239));
   MUX2_X1 i_132_0_721 (.A(\o_buffer[13] [14]), .B(i_mem_data[14]), .S(n_106), 
      .Z(n_132_238));
   MUX2_X1 i_132_0_722 (.A(\o_buffer[13] [13]), .B(i_mem_data[13]), .S(n_106), 
      .Z(n_132_237));
   MUX2_X1 i_132_0_723 (.A(\o_buffer[13] [12]), .B(i_mem_data[12]), .S(n_106), 
      .Z(n_132_236));
   MUX2_X1 i_132_0_724 (.A(\o_buffer[13] [11]), .B(i_mem_data[11]), .S(n_106), 
      .Z(n_132_235));
   MUX2_X1 i_132_0_725 (.A(\o_buffer[13] [10]), .B(i_mem_data[10]), .S(n_106), 
      .Z(n_132_234));
   MUX2_X1 i_132_0_726 (.A(\o_buffer[13] [9]), .B(i_mem_data[9]), .S(n_106), 
      .Z(n_132_233));
   MUX2_X1 i_132_0_727 (.A(\o_buffer[13] [8]), .B(i_mem_data[8]), .S(n_106), 
      .Z(n_132_232));
   MUX2_X1 i_132_0_728 (.A(\o_buffer[13] [7]), .B(i_mem_data[7]), .S(n_106), 
      .Z(n_132_231));
   MUX2_X1 i_132_0_729 (.A(\o_buffer[13] [6]), .B(i_mem_data[6]), .S(n_106), 
      .Z(n_132_230));
   MUX2_X1 i_132_0_730 (.A(\o_buffer[13] [5]), .B(i_mem_data[5]), .S(n_106), 
      .Z(n_132_229));
   MUX2_X1 i_132_0_731 (.A(\o_buffer[13] [4]), .B(i_mem_data[4]), .S(n_106), 
      .Z(n_132_228));
   MUX2_X1 i_132_0_732 (.A(\o_buffer[13] [3]), .B(i_mem_data[3]), .S(n_106), 
      .Z(n_132_227));
   MUX2_X1 i_132_0_733 (.A(\o_buffer[13] [2]), .B(i_mem_data[2]), .S(n_106), 
      .Z(n_132_226));
   MUX2_X1 i_132_0_734 (.A(\o_buffer[13] [1]), .B(i_mem_data[1]), .S(n_106), 
      .Z(n_132_225));
   MUX2_X1 i_132_0_735 (.A(\o_buffer[13] [0]), .B(i_mem_data[0]), .S(n_106), 
      .Z(n_132_224));
   MUX2_X1 i_132_0_736 (.A(\o_buffer[12] [15]), .B(i_mem_data[15]), .S(n_107), 
      .Z(n_132_223));
   MUX2_X1 i_132_0_737 (.A(\o_buffer[12] [14]), .B(i_mem_data[14]), .S(n_107), 
      .Z(n_132_222));
   MUX2_X1 i_132_0_738 (.A(\o_buffer[12] [13]), .B(i_mem_data[13]), .S(n_107), 
      .Z(n_132_221));
   MUX2_X1 i_132_0_739 (.A(\o_buffer[12] [12]), .B(i_mem_data[12]), .S(n_107), 
      .Z(n_132_220));
   MUX2_X1 i_132_0_740 (.A(\o_buffer[12] [11]), .B(i_mem_data[11]), .S(n_107), 
      .Z(n_132_219));
   MUX2_X1 i_132_0_741 (.A(\o_buffer[12] [10]), .B(i_mem_data[10]), .S(n_107), 
      .Z(n_132_218));
   MUX2_X1 i_132_0_742 (.A(\o_buffer[12] [9]), .B(i_mem_data[9]), .S(n_107), 
      .Z(n_132_217));
   MUX2_X1 i_132_0_743 (.A(\o_buffer[12] [8]), .B(i_mem_data[8]), .S(n_107), 
      .Z(n_132_216));
   MUX2_X1 i_132_0_744 (.A(\o_buffer[12] [7]), .B(i_mem_data[7]), .S(n_107), 
      .Z(n_132_215));
   MUX2_X1 i_132_0_745 (.A(\o_buffer[12] [6]), .B(i_mem_data[6]), .S(n_107), 
      .Z(n_132_214));
   MUX2_X1 i_132_0_746 (.A(\o_buffer[12] [5]), .B(i_mem_data[5]), .S(n_107), 
      .Z(n_132_213));
   MUX2_X1 i_132_0_747 (.A(\o_buffer[12] [4]), .B(i_mem_data[4]), .S(n_107), 
      .Z(n_132_212));
   MUX2_X1 i_132_0_748 (.A(\o_buffer[12] [3]), .B(i_mem_data[3]), .S(n_107), 
      .Z(n_132_211));
   MUX2_X1 i_132_0_749 (.A(\o_buffer[12] [2]), .B(i_mem_data[2]), .S(n_107), 
      .Z(n_132_210));
   MUX2_X1 i_132_0_750 (.A(\o_buffer[12] [1]), .B(i_mem_data[1]), .S(n_107), 
      .Z(n_132_209));
   MUX2_X1 i_132_0_751 (.A(\o_buffer[12] [0]), .B(i_mem_data[0]), .S(n_107), 
      .Z(n_132_208));
   MUX2_X1 i_132_0_752 (.A(\o_buffer[11] [15]), .B(i_mem_data[15]), .S(n_108), 
      .Z(n_132_207));
   MUX2_X1 i_132_0_753 (.A(\o_buffer[11] [14]), .B(i_mem_data[14]), .S(n_108), 
      .Z(n_132_206));
   MUX2_X1 i_132_0_754 (.A(\o_buffer[11] [13]), .B(i_mem_data[13]), .S(n_108), 
      .Z(n_132_205));
   MUX2_X1 i_132_0_755 (.A(\o_buffer[11] [12]), .B(i_mem_data[12]), .S(n_108), 
      .Z(n_132_204));
   MUX2_X1 i_132_0_756 (.A(\o_buffer[11] [11]), .B(i_mem_data[11]), .S(n_108), 
      .Z(n_132_203));
   MUX2_X1 i_132_0_757 (.A(\o_buffer[11] [10]), .B(i_mem_data[10]), .S(n_108), 
      .Z(n_132_202));
   MUX2_X1 i_132_0_758 (.A(\o_buffer[11] [9]), .B(i_mem_data[9]), .S(n_108), 
      .Z(n_132_201));
   MUX2_X1 i_132_0_759 (.A(\o_buffer[11] [8]), .B(i_mem_data[8]), .S(n_108), 
      .Z(n_132_200));
   MUX2_X1 i_132_0_760 (.A(\o_buffer[11] [7]), .B(i_mem_data[7]), .S(n_108), 
      .Z(n_132_199));
   MUX2_X1 i_132_0_761 (.A(\o_buffer[11] [6]), .B(i_mem_data[6]), .S(n_108), 
      .Z(n_132_198));
   MUX2_X1 i_132_0_762 (.A(\o_buffer[11] [5]), .B(i_mem_data[5]), .S(n_108), 
      .Z(n_132_197));
   MUX2_X1 i_132_0_763 (.A(\o_buffer[11] [4]), .B(i_mem_data[4]), .S(n_108), 
      .Z(n_132_196));
   MUX2_X1 i_132_0_764 (.A(\o_buffer[11] [3]), .B(i_mem_data[3]), .S(n_108), 
      .Z(n_132_195));
   MUX2_X1 i_132_0_765 (.A(\o_buffer[11] [2]), .B(i_mem_data[2]), .S(n_108), 
      .Z(n_132_194));
   MUX2_X1 i_132_0_766 (.A(\o_buffer[11] [1]), .B(i_mem_data[1]), .S(n_108), 
      .Z(n_132_193));
   MUX2_X1 i_132_0_767 (.A(\o_buffer[11] [0]), .B(i_mem_data[0]), .S(n_108), 
      .Z(n_132_192));
   MUX2_X1 i_132_0_768 (.A(\o_buffer[10] [15]), .B(i_mem_data[15]), .S(n_109), 
      .Z(n_132_191));
   MUX2_X1 i_132_0_769 (.A(\o_buffer[10] [14]), .B(i_mem_data[14]), .S(n_109), 
      .Z(n_132_190));
   MUX2_X1 i_132_0_770 (.A(\o_buffer[10] [13]), .B(i_mem_data[13]), .S(n_109), 
      .Z(n_132_189));
   MUX2_X1 i_132_0_771 (.A(\o_buffer[10] [12]), .B(i_mem_data[12]), .S(n_109), 
      .Z(n_132_188));
   MUX2_X1 i_132_0_772 (.A(\o_buffer[10] [11]), .B(i_mem_data[11]), .S(n_109), 
      .Z(n_132_187));
   MUX2_X1 i_132_0_773 (.A(\o_buffer[10] [10]), .B(i_mem_data[10]), .S(n_109), 
      .Z(n_132_186));
   MUX2_X1 i_132_0_774 (.A(\o_buffer[10] [9]), .B(i_mem_data[9]), .S(n_109), 
      .Z(n_132_185));
   MUX2_X1 i_132_0_775 (.A(\o_buffer[10] [8]), .B(i_mem_data[8]), .S(n_109), 
      .Z(n_132_184));
   MUX2_X1 i_132_0_776 (.A(\o_buffer[10] [7]), .B(i_mem_data[7]), .S(n_109), 
      .Z(n_132_183));
   MUX2_X1 i_132_0_777 (.A(\o_buffer[10] [6]), .B(i_mem_data[6]), .S(n_109), 
      .Z(n_132_182));
   MUX2_X1 i_132_0_778 (.A(\o_buffer[10] [5]), .B(i_mem_data[5]), .S(n_109), 
      .Z(n_132_181));
   MUX2_X1 i_132_0_779 (.A(\o_buffer[10] [4]), .B(i_mem_data[4]), .S(n_109), 
      .Z(n_132_180));
   MUX2_X1 i_132_0_780 (.A(\o_buffer[10] [3]), .B(i_mem_data[3]), .S(n_109), 
      .Z(n_132_179));
   MUX2_X1 i_132_0_781 (.A(\o_buffer[10] [2]), .B(i_mem_data[2]), .S(n_109), 
      .Z(n_132_178));
   MUX2_X1 i_132_0_782 (.A(\o_buffer[10] [1]), .B(i_mem_data[1]), .S(n_109), 
      .Z(n_132_177));
   MUX2_X1 i_132_0_783 (.A(\o_buffer[10] [0]), .B(i_mem_data[0]), .S(n_109), 
      .Z(n_132_176));
   MUX2_X1 i_132_0_784 (.A(\o_buffer[9] [15]), .B(i_mem_data[15]), .S(n_110), 
      .Z(n_132_175));
   MUX2_X1 i_132_0_785 (.A(\o_buffer[9] [14]), .B(i_mem_data[14]), .S(n_110), 
      .Z(n_132_174));
   MUX2_X1 i_132_0_786 (.A(\o_buffer[9] [13]), .B(i_mem_data[13]), .S(n_110), 
      .Z(n_132_173));
   MUX2_X1 i_132_0_787 (.A(\o_buffer[9] [12]), .B(i_mem_data[12]), .S(n_110), 
      .Z(n_132_172));
   MUX2_X1 i_132_0_788 (.A(\o_buffer[9] [11]), .B(i_mem_data[11]), .S(n_110), 
      .Z(n_132_171));
   MUX2_X1 i_132_0_789 (.A(\o_buffer[9] [10]), .B(i_mem_data[10]), .S(n_110), 
      .Z(n_132_170));
   MUX2_X1 i_132_0_790 (.A(\o_buffer[9] [9]), .B(i_mem_data[9]), .S(n_110), 
      .Z(n_132_169));
   MUX2_X1 i_132_0_791 (.A(\o_buffer[9] [8]), .B(i_mem_data[8]), .S(n_110), 
      .Z(n_132_168));
   MUX2_X1 i_132_0_792 (.A(\o_buffer[9] [7]), .B(i_mem_data[7]), .S(n_110), 
      .Z(n_132_167));
   MUX2_X1 i_132_0_793 (.A(\o_buffer[9] [6]), .B(i_mem_data[6]), .S(n_110), 
      .Z(n_132_166));
   MUX2_X1 i_132_0_794 (.A(\o_buffer[9] [5]), .B(i_mem_data[5]), .S(n_110), 
      .Z(n_132_165));
   MUX2_X1 i_132_0_795 (.A(\o_buffer[9] [4]), .B(i_mem_data[4]), .S(n_110), 
      .Z(n_132_164));
   MUX2_X1 i_132_0_796 (.A(\o_buffer[9] [3]), .B(i_mem_data[3]), .S(n_110), 
      .Z(n_132_163));
   MUX2_X1 i_132_0_797 (.A(\o_buffer[9] [2]), .B(i_mem_data[2]), .S(n_110), 
      .Z(n_132_162));
   MUX2_X1 i_132_0_798 (.A(\o_buffer[9] [1]), .B(i_mem_data[1]), .S(n_110), 
      .Z(n_132_161));
   MUX2_X1 i_132_0_799 (.A(\o_buffer[9] [0]), .B(i_mem_data[0]), .S(n_110), 
      .Z(n_132_160));
   MUX2_X1 i_132_0_800 (.A(\o_buffer[8] [15]), .B(i_mem_data[15]), .S(n_111), 
      .Z(n_132_159));
   MUX2_X1 i_132_0_801 (.A(\o_buffer[8] [14]), .B(i_mem_data[14]), .S(n_111), 
      .Z(n_132_158));
   MUX2_X1 i_132_0_802 (.A(\o_buffer[8] [13]), .B(i_mem_data[13]), .S(n_111), 
      .Z(n_132_157));
   MUX2_X1 i_132_0_803 (.A(\o_buffer[8] [12]), .B(i_mem_data[12]), .S(n_111), 
      .Z(n_132_156));
   MUX2_X1 i_132_0_804 (.A(\o_buffer[8] [11]), .B(i_mem_data[11]), .S(n_111), 
      .Z(n_132_155));
   MUX2_X1 i_132_0_805 (.A(\o_buffer[8] [10]), .B(i_mem_data[10]), .S(n_111), 
      .Z(n_132_154));
   MUX2_X1 i_132_0_806 (.A(\o_buffer[8] [9]), .B(i_mem_data[9]), .S(n_111), 
      .Z(n_132_153));
   MUX2_X1 i_132_0_807 (.A(\o_buffer[8] [8]), .B(i_mem_data[8]), .S(n_111), 
      .Z(n_132_152));
   MUX2_X1 i_132_0_808 (.A(\o_buffer[8] [7]), .B(i_mem_data[7]), .S(n_111), 
      .Z(n_132_151));
   MUX2_X1 i_132_0_809 (.A(\o_buffer[8] [6]), .B(i_mem_data[6]), .S(n_111), 
      .Z(n_132_150));
   MUX2_X1 i_132_0_810 (.A(\o_buffer[8] [5]), .B(i_mem_data[5]), .S(n_111), 
      .Z(n_132_149));
   MUX2_X1 i_132_0_811 (.A(\o_buffer[8] [4]), .B(i_mem_data[4]), .S(n_111), 
      .Z(n_132_148));
   MUX2_X1 i_132_0_812 (.A(\o_buffer[8] [3]), .B(i_mem_data[3]), .S(n_111), 
      .Z(n_132_147));
   MUX2_X1 i_132_0_813 (.A(\o_buffer[8] [2]), .B(i_mem_data[2]), .S(n_111), 
      .Z(n_132_146));
   MUX2_X1 i_132_0_814 (.A(\o_buffer[8] [1]), .B(i_mem_data[1]), .S(n_111), 
      .Z(n_132_145));
   MUX2_X1 i_132_0_815 (.A(\o_buffer[8] [0]), .B(i_mem_data[0]), .S(n_111), 
      .Z(n_132_144));
   MUX2_X1 i_132_0_816 (.A(\o_buffer[7] [15]), .B(i_mem_data[15]), .S(n_112), 
      .Z(n_132_143));
   MUX2_X1 i_132_0_817 (.A(\o_buffer[7] [14]), .B(i_mem_data[14]), .S(n_112), 
      .Z(n_132_142));
   MUX2_X1 i_132_0_818 (.A(\o_buffer[7] [13]), .B(i_mem_data[13]), .S(n_112), 
      .Z(n_132_141));
   MUX2_X1 i_132_0_819 (.A(\o_buffer[7] [12]), .B(i_mem_data[12]), .S(n_112), 
      .Z(n_132_140));
   MUX2_X1 i_132_0_820 (.A(\o_buffer[7] [11]), .B(i_mem_data[11]), .S(n_112), 
      .Z(n_132_139));
   MUX2_X1 i_132_0_821 (.A(\o_buffer[7] [10]), .B(i_mem_data[10]), .S(n_112), 
      .Z(n_132_138));
   MUX2_X1 i_132_0_822 (.A(\o_buffer[7] [9]), .B(i_mem_data[9]), .S(n_112), 
      .Z(n_132_137));
   MUX2_X1 i_132_0_823 (.A(\o_buffer[7] [8]), .B(i_mem_data[8]), .S(n_112), 
      .Z(n_132_136));
   MUX2_X1 i_132_0_824 (.A(\o_buffer[7] [7]), .B(i_mem_data[7]), .S(n_112), 
      .Z(n_132_135));
   MUX2_X1 i_132_0_825 (.A(\o_buffer[7] [6]), .B(i_mem_data[6]), .S(n_112), 
      .Z(n_132_134));
   MUX2_X1 i_132_0_826 (.A(\o_buffer[7] [5]), .B(i_mem_data[5]), .S(n_112), 
      .Z(n_132_133));
   MUX2_X1 i_132_0_827 (.A(\o_buffer[7] [4]), .B(i_mem_data[4]), .S(n_112), 
      .Z(n_132_132));
   MUX2_X1 i_132_0_828 (.A(\o_buffer[7] [3]), .B(i_mem_data[3]), .S(n_112), 
      .Z(n_132_131));
   MUX2_X1 i_132_0_829 (.A(\o_buffer[7] [2]), .B(i_mem_data[2]), .S(n_112), 
      .Z(n_132_130));
   MUX2_X1 i_132_0_830 (.A(\o_buffer[7] [1]), .B(i_mem_data[1]), .S(n_112), 
      .Z(n_132_129));
   MUX2_X1 i_132_0_831 (.A(\o_buffer[7] [0]), .B(i_mem_data[0]), .S(n_112), 
      .Z(n_132_128));
   MUX2_X1 i_132_0_832 (.A(\o_buffer[6] [15]), .B(i_mem_data[15]), .S(n_113), 
      .Z(n_132_127));
   MUX2_X1 i_132_0_833 (.A(\o_buffer[6] [14]), .B(i_mem_data[14]), .S(n_113), 
      .Z(n_132_126));
   MUX2_X1 i_132_0_834 (.A(\o_buffer[6] [13]), .B(i_mem_data[13]), .S(n_113), 
      .Z(n_132_125));
   MUX2_X1 i_132_0_835 (.A(\o_buffer[6] [12]), .B(i_mem_data[12]), .S(n_113), 
      .Z(n_132_124));
   MUX2_X1 i_132_0_836 (.A(\o_buffer[6] [11]), .B(i_mem_data[11]), .S(n_113), 
      .Z(n_132_123));
   MUX2_X1 i_132_0_837 (.A(\o_buffer[6] [10]), .B(i_mem_data[10]), .S(n_113), 
      .Z(n_132_122));
   MUX2_X1 i_132_0_838 (.A(\o_buffer[6] [9]), .B(i_mem_data[9]), .S(n_113), 
      .Z(n_132_121));
   MUX2_X1 i_132_0_839 (.A(\o_buffer[6] [8]), .B(i_mem_data[8]), .S(n_113), 
      .Z(n_132_120));
   MUX2_X1 i_132_0_840 (.A(\o_buffer[6] [7]), .B(i_mem_data[7]), .S(n_113), 
      .Z(n_132_119));
   MUX2_X1 i_132_0_841 (.A(\o_buffer[6] [6]), .B(i_mem_data[6]), .S(n_113), 
      .Z(n_132_118));
   MUX2_X1 i_132_0_842 (.A(\o_buffer[6] [5]), .B(i_mem_data[5]), .S(n_113), 
      .Z(n_132_117));
   MUX2_X1 i_132_0_843 (.A(\o_buffer[6] [4]), .B(i_mem_data[4]), .S(n_113), 
      .Z(n_132_116));
   MUX2_X1 i_132_0_844 (.A(\o_buffer[6] [3]), .B(i_mem_data[3]), .S(n_113), 
      .Z(n_132_115));
   MUX2_X1 i_132_0_845 (.A(\o_buffer[6] [2]), .B(i_mem_data[2]), .S(n_113), 
      .Z(n_132_114));
   MUX2_X1 i_132_0_846 (.A(\o_buffer[6] [1]), .B(i_mem_data[1]), .S(n_113), 
      .Z(n_132_113));
   MUX2_X1 i_132_0_847 (.A(\o_buffer[6] [0]), .B(i_mem_data[0]), .S(n_113), 
      .Z(n_132_112));
   MUX2_X1 i_132_0_848 (.A(\o_buffer[5] [15]), .B(i_mem_data[15]), .S(n_114), 
      .Z(n_132_111));
   MUX2_X1 i_132_0_849 (.A(\o_buffer[5] [14]), .B(i_mem_data[14]), .S(n_114), 
      .Z(n_132_110));
   MUX2_X1 i_132_0_850 (.A(\o_buffer[5] [13]), .B(i_mem_data[13]), .S(n_114), 
      .Z(n_132_109));
   MUX2_X1 i_132_0_851 (.A(\o_buffer[5] [12]), .B(i_mem_data[12]), .S(n_114), 
      .Z(n_132_108));
   MUX2_X1 i_132_0_852 (.A(\o_buffer[5] [11]), .B(i_mem_data[11]), .S(n_114), 
      .Z(n_132_107));
   MUX2_X1 i_132_0_853 (.A(\o_buffer[5] [10]), .B(i_mem_data[10]), .S(n_114), 
      .Z(n_132_106));
   MUX2_X1 i_132_0_854 (.A(\o_buffer[5] [9]), .B(i_mem_data[9]), .S(n_114), 
      .Z(n_132_105));
   MUX2_X1 i_132_0_855 (.A(\o_buffer[5] [8]), .B(i_mem_data[8]), .S(n_114), 
      .Z(n_132_104));
   MUX2_X1 i_132_0_856 (.A(\o_buffer[5] [7]), .B(i_mem_data[7]), .S(n_114), 
      .Z(n_132_103));
   MUX2_X1 i_132_0_857 (.A(\o_buffer[5] [6]), .B(i_mem_data[6]), .S(n_114), 
      .Z(n_132_102));
   MUX2_X1 i_132_0_858 (.A(\o_buffer[5] [5]), .B(i_mem_data[5]), .S(n_114), 
      .Z(n_132_101));
   MUX2_X1 i_132_0_859 (.A(\o_buffer[5] [4]), .B(i_mem_data[4]), .S(n_114), 
      .Z(n_132_100));
   MUX2_X1 i_132_0_860 (.A(\o_buffer[5] [3]), .B(i_mem_data[3]), .S(n_114), 
      .Z(n_132_99));
   MUX2_X1 i_132_0_861 (.A(\o_buffer[5] [2]), .B(i_mem_data[2]), .S(n_114), 
      .Z(n_132_98));
   MUX2_X1 i_132_0_862 (.A(\o_buffer[5] [1]), .B(i_mem_data[1]), .S(n_114), 
      .Z(n_132_97));
   MUX2_X1 i_132_0_863 (.A(\o_buffer[5] [0]), .B(i_mem_data[0]), .S(n_114), 
      .Z(n_132_96));
   MUX2_X1 i_132_0_864 (.A(\o_buffer[4] [15]), .B(i_mem_data[15]), .S(n_115), 
      .Z(n_132_95));
   MUX2_X1 i_132_0_865 (.A(\o_buffer[4] [14]), .B(i_mem_data[14]), .S(n_115), 
      .Z(n_132_94));
   MUX2_X1 i_132_0_866 (.A(\o_buffer[4] [13]), .B(i_mem_data[13]), .S(n_115), 
      .Z(n_132_93));
   MUX2_X1 i_132_0_867 (.A(\o_buffer[4] [12]), .B(i_mem_data[12]), .S(n_115), 
      .Z(n_132_92));
   MUX2_X1 i_132_0_868 (.A(\o_buffer[4] [11]), .B(i_mem_data[11]), .S(n_115), 
      .Z(n_132_91));
   MUX2_X1 i_132_0_869 (.A(\o_buffer[4] [10]), .B(i_mem_data[10]), .S(n_115), 
      .Z(n_132_90));
   MUX2_X1 i_132_0_870 (.A(\o_buffer[4] [9]), .B(i_mem_data[9]), .S(n_115), 
      .Z(n_132_89));
   MUX2_X1 i_132_0_871 (.A(\o_buffer[4] [8]), .B(i_mem_data[8]), .S(n_115), 
      .Z(n_132_88));
   MUX2_X1 i_132_0_872 (.A(\o_buffer[4] [7]), .B(i_mem_data[7]), .S(n_115), 
      .Z(n_132_87));
   MUX2_X1 i_132_0_873 (.A(\o_buffer[4] [6]), .B(i_mem_data[6]), .S(n_115), 
      .Z(n_132_86));
   MUX2_X1 i_132_0_874 (.A(\o_buffer[4] [5]), .B(i_mem_data[5]), .S(n_115), 
      .Z(n_132_85));
   MUX2_X1 i_132_0_875 (.A(\o_buffer[4] [4]), .B(i_mem_data[4]), .S(n_115), 
      .Z(n_132_84));
   MUX2_X1 i_132_0_876 (.A(\o_buffer[4] [3]), .B(i_mem_data[3]), .S(n_115), 
      .Z(n_132_83));
   MUX2_X1 i_132_0_877 (.A(\o_buffer[4] [2]), .B(i_mem_data[2]), .S(n_115), 
      .Z(n_132_82));
   MUX2_X1 i_132_0_878 (.A(\o_buffer[4] [1]), .B(i_mem_data[1]), .S(n_115), 
      .Z(n_132_81));
   MUX2_X1 i_132_0_879 (.A(\o_buffer[4] [0]), .B(i_mem_data[0]), .S(n_115), 
      .Z(n_132_80));
   MUX2_X1 i_132_0_880 (.A(\o_buffer[3] [15]), .B(i_mem_data[15]), .S(n_116), 
      .Z(n_132_79));
   MUX2_X1 i_132_0_881 (.A(\o_buffer[3] [14]), .B(i_mem_data[14]), .S(n_116), 
      .Z(n_132_78));
   MUX2_X1 i_132_0_882 (.A(\o_buffer[3] [13]), .B(i_mem_data[13]), .S(n_116), 
      .Z(n_132_77));
   MUX2_X1 i_132_0_883 (.A(\o_buffer[3] [12]), .B(i_mem_data[12]), .S(n_116), 
      .Z(n_132_76));
   MUX2_X1 i_132_0_884 (.A(\o_buffer[3] [11]), .B(i_mem_data[11]), .S(n_116), 
      .Z(n_132_75));
   MUX2_X1 i_132_0_885 (.A(\o_buffer[3] [10]), .B(i_mem_data[10]), .S(n_116), 
      .Z(n_132_74));
   MUX2_X1 i_132_0_886 (.A(\o_buffer[3] [9]), .B(i_mem_data[9]), .S(n_116), 
      .Z(n_132_73));
   MUX2_X1 i_132_0_887 (.A(\o_buffer[3] [8]), .B(i_mem_data[8]), .S(n_116), 
      .Z(n_132_72));
   MUX2_X1 i_132_0_888 (.A(\o_buffer[3] [7]), .B(i_mem_data[7]), .S(n_116), 
      .Z(n_132_71));
   MUX2_X1 i_132_0_889 (.A(\o_buffer[3] [6]), .B(i_mem_data[6]), .S(n_116), 
      .Z(n_132_70));
   MUX2_X1 i_132_0_890 (.A(\o_buffer[3] [5]), .B(i_mem_data[5]), .S(n_116), 
      .Z(n_132_69));
   MUX2_X1 i_132_0_891 (.A(\o_buffer[3] [4]), .B(i_mem_data[4]), .S(n_116), 
      .Z(n_132_68));
   MUX2_X1 i_132_0_892 (.A(\o_buffer[3] [3]), .B(i_mem_data[3]), .S(n_116), 
      .Z(n_132_67));
   MUX2_X1 i_132_0_893 (.A(\o_buffer[3] [2]), .B(i_mem_data[2]), .S(n_116), 
      .Z(n_132_66));
   MUX2_X1 i_132_0_894 (.A(\o_buffer[3] [1]), .B(i_mem_data[1]), .S(n_116), 
      .Z(n_132_65));
   MUX2_X1 i_132_0_895 (.A(\o_buffer[3] [0]), .B(i_mem_data[0]), .S(n_116), 
      .Z(n_132_64));
   MUX2_X1 i_132_0_896 (.A(\o_buffer[2] [15]), .B(i_mem_data[15]), .S(n_117), 
      .Z(n_132_63));
   MUX2_X1 i_132_0_897 (.A(\o_buffer[2] [14]), .B(i_mem_data[14]), .S(n_117), 
      .Z(n_132_62));
   MUX2_X1 i_132_0_898 (.A(\o_buffer[2] [13]), .B(i_mem_data[13]), .S(n_117), 
      .Z(n_132_61));
   MUX2_X1 i_132_0_899 (.A(\o_buffer[2] [12]), .B(i_mem_data[12]), .S(n_117), 
      .Z(n_132_60));
   MUX2_X1 i_132_0_900 (.A(\o_buffer[2] [11]), .B(i_mem_data[11]), .S(n_117), 
      .Z(n_132_59));
   MUX2_X1 i_132_0_901 (.A(\o_buffer[2] [10]), .B(i_mem_data[10]), .S(n_117), 
      .Z(n_132_58));
   MUX2_X1 i_132_0_902 (.A(\o_buffer[2] [9]), .B(i_mem_data[9]), .S(n_117), 
      .Z(n_132_57));
   MUX2_X1 i_132_0_903 (.A(\o_buffer[2] [8]), .B(i_mem_data[8]), .S(n_117), 
      .Z(n_132_56));
   MUX2_X1 i_132_0_904 (.A(\o_buffer[2] [7]), .B(i_mem_data[7]), .S(n_117), 
      .Z(n_132_55));
   MUX2_X1 i_132_0_905 (.A(\o_buffer[2] [6]), .B(i_mem_data[6]), .S(n_117), 
      .Z(n_132_54));
   MUX2_X1 i_132_0_906 (.A(\o_buffer[2] [5]), .B(i_mem_data[5]), .S(n_117), 
      .Z(n_132_53));
   MUX2_X1 i_132_0_907 (.A(\o_buffer[2] [4]), .B(i_mem_data[4]), .S(n_117), 
      .Z(n_132_52));
   MUX2_X1 i_132_0_908 (.A(\o_buffer[2] [3]), .B(i_mem_data[3]), .S(n_117), 
      .Z(n_132_51));
   MUX2_X1 i_132_0_909 (.A(\o_buffer[2] [2]), .B(i_mem_data[2]), .S(n_117), 
      .Z(n_132_50));
   MUX2_X1 i_132_0_910 (.A(\o_buffer[2] [1]), .B(i_mem_data[1]), .S(n_117), 
      .Z(n_132_49));
   MUX2_X1 i_132_0_911 (.A(\o_buffer[2] [0]), .B(i_mem_data[0]), .S(n_117), 
      .Z(n_132_48));
   MUX2_X1 i_132_0_912 (.A(\o_buffer[1] [15]), .B(i_mem_data[15]), .S(n_118), 
      .Z(n_132_47));
   MUX2_X1 i_132_0_913 (.A(\o_buffer[1] [14]), .B(i_mem_data[14]), .S(n_118), 
      .Z(n_132_46));
   MUX2_X1 i_132_0_914 (.A(\o_buffer[1] [13]), .B(i_mem_data[13]), .S(n_118), 
      .Z(n_132_45));
   MUX2_X1 i_132_0_915 (.A(\o_buffer[1] [12]), .B(i_mem_data[12]), .S(n_118), 
      .Z(n_132_44));
   MUX2_X1 i_132_0_916 (.A(\o_buffer[1] [11]), .B(i_mem_data[11]), .S(n_118), 
      .Z(n_132_43));
   MUX2_X1 i_132_0_917 (.A(\o_buffer[1] [10]), .B(i_mem_data[10]), .S(n_118), 
      .Z(n_132_42));
   MUX2_X1 i_132_0_918 (.A(\o_buffer[1] [9]), .B(i_mem_data[9]), .S(n_118), 
      .Z(n_132_41));
   MUX2_X1 i_132_0_919 (.A(\o_buffer[1] [8]), .B(i_mem_data[8]), .S(n_118), 
      .Z(n_132_40));
   MUX2_X1 i_132_0_920 (.A(\o_buffer[1] [7]), .B(i_mem_data[7]), .S(n_118), 
      .Z(n_132_39));
   MUX2_X1 i_132_0_921 (.A(\o_buffer[1] [6]), .B(i_mem_data[6]), .S(n_118), 
      .Z(n_132_38));
   MUX2_X1 i_132_0_922 (.A(\o_buffer[1] [5]), .B(i_mem_data[5]), .S(n_118), 
      .Z(n_132_37));
   MUX2_X1 i_132_0_923 (.A(\o_buffer[1] [4]), .B(i_mem_data[4]), .S(n_118), 
      .Z(n_132_36));
   MUX2_X1 i_132_0_924 (.A(\o_buffer[1] [3]), .B(i_mem_data[3]), .S(n_118), 
      .Z(n_132_35));
   MUX2_X1 i_132_0_925 (.A(\o_buffer[1] [2]), .B(i_mem_data[2]), .S(n_118), 
      .Z(n_132_34));
   MUX2_X1 i_132_0_926 (.A(\o_buffer[1] [1]), .B(i_mem_data[1]), .S(n_118), 
      .Z(n_132_33));
   MUX2_X1 i_132_0_927 (.A(\o_buffer[1] [0]), .B(i_mem_data[0]), .S(n_118), 
      .Z(n_132_32));
   MUX2_X1 i_132_0_928 (.A(\o_buffer[0] [15]), .B(i_mem_data[15]), .S(n_119), 
      .Z(n_132_31));
   MUX2_X1 i_132_0_929 (.A(\o_buffer[0] [14]), .B(i_mem_data[14]), .S(n_119), 
      .Z(n_132_30));
   MUX2_X1 i_132_0_930 (.A(\o_buffer[0] [13]), .B(i_mem_data[13]), .S(n_119), 
      .Z(n_132_29));
   MUX2_X1 i_132_0_931 (.A(\o_buffer[0] [12]), .B(i_mem_data[12]), .S(n_119), 
      .Z(n_132_28));
   MUX2_X1 i_132_0_932 (.A(\o_buffer[0] [11]), .B(i_mem_data[11]), .S(n_119), 
      .Z(n_132_27));
   MUX2_X1 i_132_0_933 (.A(\o_buffer[0] [10]), .B(i_mem_data[10]), .S(n_119), 
      .Z(n_132_26));
   MUX2_X1 i_132_0_934 (.A(\o_buffer[0] [9]), .B(i_mem_data[9]), .S(n_119), 
      .Z(n_132_25));
   MUX2_X1 i_132_0_935 (.A(\o_buffer[0] [8]), .B(i_mem_data[8]), .S(n_119), 
      .Z(n_132_24));
   MUX2_X1 i_132_0_936 (.A(\o_buffer[0] [7]), .B(i_mem_data[7]), .S(n_119), 
      .Z(n_132_23));
   MUX2_X1 i_132_0_937 (.A(\o_buffer[0] [6]), .B(i_mem_data[6]), .S(n_119), 
      .Z(n_132_22));
   MUX2_X1 i_132_0_938 (.A(\o_buffer[0] [5]), .B(i_mem_data[5]), .S(n_119), 
      .Z(n_132_21));
   MUX2_X1 i_132_0_939 (.A(\o_buffer[0] [4]), .B(i_mem_data[4]), .S(n_119), 
      .Z(n_132_20));
   MUX2_X1 i_132_0_940 (.A(\o_buffer[0] [3]), .B(i_mem_data[3]), .S(n_119), 
      .Z(n_132_19));
   MUX2_X1 i_132_0_941 (.A(\o_buffer[0] [2]), .B(i_mem_data[2]), .S(n_119), 
      .Z(n_132_18));
   MUX2_X1 i_132_0_942 (.A(\o_buffer[0] [1]), .B(i_mem_data[1]), .S(n_119), 
      .Z(n_132_17));
   MUX2_X1 i_132_0_943 (.A(\o_buffer[0] [0]), .B(i_mem_data[0]), .S(n_119), 
      .Z(n_132_16));
   MUX2_X1 i_132_0_944 (.A(\o_buffer[119] [15]), .B(i_mem_data[15]), .S(n_0), 
      .Z(n_132_15));
   MUX2_X1 i_132_0_945 (.A(\o_buffer[119] [14]), .B(i_mem_data[14]), .S(n_0), 
      .Z(n_132_14));
   MUX2_X1 i_132_0_946 (.A(\o_buffer[119] [13]), .B(i_mem_data[13]), .S(n_0), 
      .Z(n_132_13));
   MUX2_X1 i_132_0_947 (.A(\o_buffer[119] [12]), .B(i_mem_data[12]), .S(n_0), 
      .Z(n_132_12));
   MUX2_X1 i_132_0_948 (.A(\o_buffer[119] [11]), .B(i_mem_data[11]), .S(n_0), 
      .Z(n_132_11));
   MUX2_X1 i_132_0_949 (.A(\o_buffer[119] [10]), .B(i_mem_data[10]), .S(n_0), 
      .Z(n_132_10));
   MUX2_X1 i_132_0_950 (.A(\o_buffer[119] [9]), .B(i_mem_data[9]), .S(n_0), 
      .Z(n_132_9));
   MUX2_X1 i_132_0_951 (.A(\o_buffer[119] [8]), .B(i_mem_data[8]), .S(n_0), 
      .Z(n_132_8));
   MUX2_X1 i_132_0_952 (.A(\o_buffer[119] [7]), .B(i_mem_data[7]), .S(n_0), 
      .Z(n_132_7));
   MUX2_X1 i_132_0_953 (.A(\o_buffer[119] [6]), .B(i_mem_data[6]), .S(n_0), 
      .Z(n_132_6));
   MUX2_X1 i_132_0_954 (.A(\o_buffer[119] [5]), .B(i_mem_data[5]), .S(n_0), 
      .Z(n_132_5));
   MUX2_X1 i_132_0_955 (.A(\o_buffer[119] [4]), .B(i_mem_data[4]), .S(n_0), 
      .Z(n_132_4));
   MUX2_X1 i_132_0_956 (.A(\o_buffer[119] [3]), .B(i_mem_data[3]), .S(n_0), 
      .Z(n_132_3));
   MUX2_X1 i_132_0_957 (.A(\o_buffer[119] [2]), .B(i_mem_data[2]), .S(n_0), 
      .Z(n_132_2));
   MUX2_X1 i_132_0_958 (.A(\o_buffer[119] [1]), .B(i_mem_data[1]), .S(n_0), 
      .Z(n_132_1));
   MUX2_X1 i_132_0_959 (.A(\o_buffer[119] [0]), .B(i_mem_data[0]), .S(n_0), 
      .Z(n_132_0));
   datapath__0_120 i_0_122 (.mem_idx({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0}), .p_0({n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, 
      n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
      n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, uc_0}));
   DFF_X1 \mem_idx_reg[31]  (.D(n_0_33), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[30]  (.D(n_0_34), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[29]  (.D(n_0_35), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[28]  (.D(n_0_36), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[27]  (.D(n_0_37), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[26]  (.D(n_0_38), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[25]  (.D(n_0_39), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[24]  (.D(n_0_40), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[23]  (.D(n_0_41), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[22]  (.D(n_0_42), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[21]  (.D(n_0_43), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[20]  (.D(n_0_44), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[19]  (.D(n_0_45), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[18]  (.D(n_0_46), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[17]  (.D(n_0_47), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[16]  (.D(n_0_48), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[15]  (.D(n_0_49), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[14]  (.D(n_0_50), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[13]  (.D(n_0_51), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[12]  (.D(n_0_52), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[11]  (.D(n_0_53), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[10]  (.D(n_0_54), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[9]  (.D(n_0_55), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[8]  (.D(n_0_56), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[7]  (.D(n_0_57), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[6]  (.D(n_0_58), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[5]  (.D(n_0_59), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[4]  (.D(n_0_60), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[3]  (.D(n_0_61), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[2]  (.D(n_0_62), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[1]  (.D(n_0_1), .CK(n_120), .Q(1'b0), .QN());
   DFF_X1 \mem_idx_reg[0]  (.D(n_0_0), .CK(n_120), .Q(1'b0), .QN());
   INV_X1 i_0_0_0 (.A(1'b0), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_1 (.A1(n_0_0_0), .A2(count[6]), .ZN(n_0_0_1));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(n_0_0_2));
   INV_X1 i_0_0_3 (.A(1'b0), .ZN(n_0_0_3));
   INV_X1 i_0_0_4 (.A(1'b0), .ZN(n_0_0_4));
   AOI221_X1 i_0_0_5 (.A(n_0_0_2), .B1(count[4]), .B2(n_0_0_3), .C1(count[5]), 
      .C2(n_0_0_4), .ZN(n_0_0_5));
   OR2_X1 i_0_0_6 (.A1(n_0_0_3), .A2(count[4]), .ZN(n_0_0_6));
   NAND2_X1 i_0_0_7 (.A1(n_0_0_6), .A2(count[3]), .ZN(n_0_0_7));
   INV_X1 i_0_0_8 (.A(1'b0), .ZN(n_0_0_8));
   INV_X1 i_0_0_9 (.A(1'b0), .ZN(n_0_0_9));
   OAI221_X1 i_0_0_10 (.A(n_0_0_6), .B1(n_0_0_8), .B2(count[2]), .C1(count[3]), 
      .C2(n_0_0_9), .ZN(n_0_0_10));
   INV_X1 i_0_0_11 (.A(count[0]), .ZN(n_0_0_11));
   OAI21_X1 i_0_0_12 (.A(1'b0), .B1(n_0_0_11), .B2(1'b0), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_13 (.A1(1'b0), .A2(1'b0), .ZN(n_0_0_13));
   AOI222_X1 i_0_0_14 (.A1(n_0_0_12), .A2(count[1]), .B1(n_0_0_13), .B2(count[0]), 
      .C1(n_0_0_8), .C2(count[2]), .ZN(n_0_0_14));
   OAI221_X1 i_0_0_15 (.A(n_0_0_5), .B1(1'b0), .B2(n_0_0_7), .C1(n_0_0_10), 
      .C2(n_0_0_14), .ZN(n_0_0_15));
   OAI22_X1 i_0_0_16 (.A1(n_0_0_4), .A2(count[5]), .B1(n_0_0_0), .B2(count[6]), 
      .ZN(n_0_0_16));
   INV_X1 i_0_0_17 (.A(count[7]), .ZN(n_0_0_17));
   AOI22_X1 i_0_0_18 (.A1(n_0_0_16), .A2(n_0_0_1), .B1(n_0_0_17), .B2(1'b0), 
      .ZN(n_0_0_18));
   INV_X1 i_0_0_19 (.A(1'b0), .ZN(n_0_0_19));
   INV_X1 i_0_0_20 (.A(1'b0), .ZN(n_0_0_20));
   AOI222_X1 i_0_0_21 (.A1(n_0_0_15), .A2(n_0_0_18), .B1(count[8]), .B2(n_0_0_19), 
      .C1(count[7]), .C2(n_0_0_20), .ZN(n_0_0_21));
   INV_X1 i_0_0_22 (.A(1'b0), .ZN(n_0_0_22));
   OAI22_X1 i_0_0_23 (.A1(n_0_0_22), .A2(count[9]), .B1(n_0_0_19), .B2(count[8]), 
      .ZN(n_0_0_23));
   INV_X1 i_0_0_24 (.A(count[9]), .ZN(n_0_0_24));
   OAI22_X1 i_0_0_25 (.A1(n_0_0_21), .A2(n_0_0_23), .B1(n_0_0_24), .B2(1'b0), 
      .ZN(n_0_0_25));
   NOR4_X1 i_0_0_26 (.A1(1'b0), .A2(1'b0), .A3(1'b0), .A4(1'b0), .ZN(n_0_0_26));
   NAND2_X1 i_0_0_27 (.A1(n_0_0_26), .A2(read), .ZN(n_0_0_27));
   OR3_X1 i_0_0_28 (.A1(n_0_0_27), .A2(1'b0), .A3(1'b0), .ZN(n_0_0_28));
   NOR4_X1 i_0_0_29 (.A1(1'b0), .A2(1'b0), .A3(1'b0), .A4(1'b0), .ZN(n_0_0_29));
   NOR4_X1 i_0_0_30 (.A1(1'b0), .A2(1'b0), .A3(1'b0), .A4(1'b0), .ZN(n_0_0_30));
   NOR4_X1 i_0_0_31 (.A1(1'b0), .A2(1'b0), .A3(1'b0), .A4(1'b0), .ZN(n_0_0_31));
   NOR3_X1 i_0_0_32 (.A1(1'b0), .A2(1'b0), .A3(1'b0), .ZN(n_0_0_32));
   NAND4_X1 i_0_0_33 (.A1(n_0_0_29), .A2(n_0_0_30), .A3(n_0_0_31), .A4(n_0_0_32), 
      .ZN(n_0_0_33));
   NOR3_X1 i_0_0_34 (.A1(n_0_0_28), .A2(1'b0), .A3(n_0_0_33), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_25), .A2(n_0_0_34), .ZN(n_0_0_35));
   INV_X1 i_0_0_36 (.A(n_0_0_35), .ZN(n_0_0_36));
   INV_X1 i_0_0_37 (.A(1'b0), .ZN(n_0_0_37));
   AOI22_X1 i_0_0_38 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_0_37), 
      .ZN(n_0_0));
   OAI22_X1 i_0_0_39 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_2), 
      .ZN(n_0_0_38));
   INV_X1 i_0_0_40 (.A(n_0_0_38), .ZN(n_0_1));
   AOI22_X1 i_0_0_41 (.A1(n_0_0_36), .A2(n_0_3), .B1(n_0_0_35), .B2(1'b0), 
      .ZN(n_0_0_39));
   INV_X1 i_0_0_42 (.A(n_0_0_39), .ZN(n_0_62));
   AOI22_X1 i_0_0_43 (.A1(n_0_0_36), .A2(n_0_4), .B1(n_0_0_35), .B2(1'b0), 
      .ZN(n_0_0_40));
   INV_X1 i_0_0_44 (.A(n_0_0_40), .ZN(n_0_61));
   AOI22_X1 i_0_0_45 (.A1(n_0_0_36), .A2(n_0_5), .B1(n_0_0_35), .B2(1'b0), 
      .ZN(n_0_0_41));
   INV_X1 i_0_0_46 (.A(n_0_0_41), .ZN(n_0_60));
   OAI22_X1 i_0_0_47 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_6), 
      .ZN(n_0_0_42));
   INV_X1 i_0_0_48 (.A(n_0_0_42), .ZN(n_0_59));
   AOI22_X1 i_0_0_49 (.A1(n_0_0_36), .A2(n_0_7), .B1(n_0_0_35), .B2(1'b0), 
      .ZN(n_0_0_43));
   INV_X1 i_0_0_50 (.A(n_0_0_43), .ZN(n_0_58));
   OAI22_X1 i_0_0_51 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_8), 
      .ZN(n_0_0_44));
   INV_X1 i_0_0_52 (.A(n_0_0_44), .ZN(n_0_57));
   OAI22_X1 i_0_0_53 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_9), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_54 (.A(n_0_0_45), .ZN(n_0_56));
   OAI22_X1 i_0_0_55 (.A1(n_0_0_36), .A2(1'b0), .B1(n_0_0_35), .B2(n_0_10), 
      .ZN(n_0_0_46));
   INV_X1 i_0_0_56 (.A(n_0_0_46), .ZN(n_0_55));
   AOI21_X1 i_0_0_57 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_11), .ZN(n_0_0_47));
   INV_X1 i_0_0_58 (.A(n_0_0_47), .ZN(n_0_54));
   AOI21_X1 i_0_0_59 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_12), .ZN(n_0_0_48));
   INV_X1 i_0_0_60 (.A(n_0_0_48), .ZN(n_0_53));
   AOI21_X1 i_0_0_61 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_13), .ZN(n_0_0_49));
   INV_X1 i_0_0_62 (.A(n_0_0_49), .ZN(n_0_52));
   AOI21_X1 i_0_0_63 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_14), .ZN(n_0_0_50));
   INV_X1 i_0_0_64 (.A(n_0_0_50), .ZN(n_0_51));
   AOI21_X1 i_0_0_65 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_15), .ZN(n_0_0_51));
   INV_X1 i_0_0_66 (.A(n_0_0_51), .ZN(n_0_50));
   AOI21_X1 i_0_0_67 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_16), .ZN(n_0_0_52));
   INV_X1 i_0_0_68 (.A(n_0_0_52), .ZN(n_0_49));
   AOI21_X1 i_0_0_69 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_17), .ZN(n_0_0_53));
   INV_X1 i_0_0_70 (.A(n_0_0_53), .ZN(n_0_48));
   AOI21_X1 i_0_0_71 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_18), .ZN(n_0_0_54));
   INV_X1 i_0_0_72 (.A(n_0_0_54), .ZN(n_0_47));
   AOI21_X1 i_0_0_73 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_19), .ZN(n_0_0_55));
   INV_X1 i_0_0_74 (.A(n_0_0_55), .ZN(n_0_46));
   AOI21_X1 i_0_0_75 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_20), .ZN(n_0_0_56));
   INV_X1 i_0_0_76 (.A(n_0_0_56), .ZN(n_0_45));
   AOI21_X1 i_0_0_77 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_21), .ZN(n_0_0_57));
   INV_X1 i_0_0_78 (.A(n_0_0_57), .ZN(n_0_44));
   AOI21_X1 i_0_0_79 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_22), .ZN(n_0_0_58));
   INV_X1 i_0_0_80 (.A(n_0_0_58), .ZN(n_0_43));
   AOI21_X1 i_0_0_81 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_23), .ZN(n_0_0_59));
   INV_X1 i_0_0_82 (.A(n_0_0_59), .ZN(n_0_42));
   AOI21_X1 i_0_0_83 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_24), .ZN(n_0_0_60));
   INV_X1 i_0_0_84 (.A(n_0_0_60), .ZN(n_0_41));
   AOI21_X1 i_0_0_85 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_25), .ZN(n_0_0_61));
   INV_X1 i_0_0_86 (.A(n_0_0_61), .ZN(n_0_40));
   AOI21_X1 i_0_0_87 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_26), .ZN(n_0_0_62));
   INV_X1 i_0_0_88 (.A(n_0_0_62), .ZN(n_0_39));
   AOI21_X1 i_0_0_89 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_27), .ZN(n_0_0_63));
   INV_X1 i_0_0_90 (.A(n_0_0_63), .ZN(n_0_38));
   AOI21_X1 i_0_0_91 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_28), .ZN(n_0_0_64));
   INV_X1 i_0_0_92 (.A(n_0_0_64), .ZN(n_0_37));
   AOI21_X1 i_0_0_93 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_29), .ZN(n_0_0_65));
   INV_X1 i_0_0_94 (.A(n_0_0_65), .ZN(n_0_36));
   AOI21_X1 i_0_0_95 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_30), .ZN(n_0_0_66));
   INV_X1 i_0_0_96 (.A(n_0_0_66), .ZN(n_0_35));
   AOI21_X1 i_0_0_97 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_31), .ZN(n_0_0_67));
   INV_X1 i_0_0_98 (.A(n_0_0_67), .ZN(n_0_34));
   AOI21_X1 i_0_0_99 (.A(1'b0), .B1(n_0_0_36), .B2(n_0_32), .ZN(n_0_0_68));
   INV_X1 i_0_0_100 (.A(n_0_0_68), .ZN(n_0_33));
   NAND4_X1 i_0_0_101 (.A1(n_0_0_36), .A2(n_0_0_19), .A3(n_0_0_20), .A4(n_0_0_22), 
      .ZN(n_0_0_69));
   NOR2_X1 i_0_0_102 (.A1(n_0_0_69), .A2(n_0_0_0), .ZN(n_0_0_70));
   NAND3_X1 i_0_0_103 (.A1(n_0_0_70), .A2(1'b0), .A3(1'b0), .ZN(n_0_0_71));
   INV_X1 i_0_0_104 (.A(1'b0), .ZN(n_0_0_72));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_37), .A2(n_0_0_72), .ZN(n_0_0_73));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_4), .A2(1'b0), .ZN(n_0_0_74));
   NAND2_X1 i_0_0_107 (.A1(n_0_0_73), .A2(n_0_0_74), .ZN(n_0_0_75));
   NOR2_X1 i_0_0_108 (.A1(n_0_0_71), .A2(n_0_0_75), .ZN(n_0));
   NOR2_X1 i_0_0_109 (.A1(n_0_0_72), .A2(1'b0), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_110 (.A1(n_0_0_74), .A2(n_0_0_76), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_111 (.A1(n_0_0_71), .A2(n_0_0_77), .ZN(n_1));
   NOR2_X1 i_0_0_112 (.A1(n_0_0_37), .A2(1'b0), .ZN(n_0_0_78));
   NAND2_X1 i_0_0_113 (.A1(n_0_0_74), .A2(n_0_0_78), .ZN(n_0_0_79));
   NOR2_X1 i_0_0_114 (.A1(n_0_0_71), .A2(n_0_0_79), .ZN(n_2));
   NAND2_X1 i_0_0_115 (.A1(n_0_0_74), .A2(n_0_0_13), .ZN(n_0_0_80));
   NOR2_X1 i_0_0_116 (.A1(n_0_0_71), .A2(n_0_0_80), .ZN(n_3));
   NAND3_X1 i_0_0_117 (.A1(n_0_0_70), .A2(1'b0), .A3(n_0_0_8), .ZN(n_0_0_81));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_81), .A2(n_0_0_75), .ZN(n_4));
   NOR2_X1 i_0_0_119 (.A1(n_0_0_81), .A2(n_0_0_77), .ZN(n_5));
   NOR2_X1 i_0_0_120 (.A1(n_0_0_81), .A2(n_0_0_79), .ZN(n_6));
   NOR2_X1 i_0_0_121 (.A1(n_0_0_81), .A2(n_0_0_80), .ZN(n_7));
   NAND3_X1 i_0_0_122 (.A1(n_0_0_70), .A2(n_0_0_3), .A3(1'b0), .ZN(n_0_0_82));
   NOR2_X1 i_0_0_123 (.A1(n_0_0_4), .A2(n_0_0_9), .ZN(n_0_0_83));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_73), .A2(n_0_0_83), .ZN(n_0_0_84));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_82), .A2(n_0_0_84), .ZN(n_8));
   NAND2_X1 i_0_0_126 (.A1(n_0_0_83), .A2(n_0_0_76), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_127 (.A1(n_0_0_82), .A2(n_0_0_85), .ZN(n_9));
   NAND2_X1 i_0_0_128 (.A1(n_0_0_83), .A2(n_0_0_78), .ZN(n_0_0_86));
   NOR2_X1 i_0_0_129 (.A1(n_0_0_82), .A2(n_0_0_86), .ZN(n_10));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_83), .A2(n_0_0_13), .ZN(n_0_0_87));
   NOR2_X1 i_0_0_131 (.A1(n_0_0_82), .A2(n_0_0_87), .ZN(n_11));
   NAND3_X1 i_0_0_132 (.A1(n_0_0_70), .A2(n_0_0_3), .A3(n_0_0_8), .ZN(n_0_0_88));
   NOR2_X1 i_0_0_133 (.A1(n_0_0_88), .A2(n_0_0_84), .ZN(n_12));
   NOR2_X1 i_0_0_134 (.A1(n_0_0_88), .A2(n_0_0_85), .ZN(n_13));
   NOR2_X1 i_0_0_135 (.A1(n_0_0_88), .A2(n_0_0_86), .ZN(n_14));
   NOR2_X1 i_0_0_136 (.A1(n_0_0_88), .A2(n_0_0_87), .ZN(n_15));
   NOR2_X1 i_0_0_137 (.A1(n_0_0_82), .A2(n_0_0_75), .ZN(n_16));
   NOR2_X1 i_0_0_138 (.A1(n_0_0_82), .A2(n_0_0_77), .ZN(n_17));
   NOR2_X1 i_0_0_139 (.A1(n_0_0_82), .A2(n_0_0_79), .ZN(n_18));
   NOR2_X1 i_0_0_140 (.A1(n_0_0_82), .A2(n_0_0_80), .ZN(n_19));
   NOR2_X1 i_0_0_141 (.A1(n_0_0_88), .A2(n_0_0_75), .ZN(n_20));
   NOR2_X1 i_0_0_142 (.A1(n_0_0_88), .A2(n_0_0_77), .ZN(n_21));
   NOR2_X1 i_0_0_143 (.A1(n_0_0_88), .A2(n_0_0_79), .ZN(n_22));
   NOR2_X1 i_0_0_144 (.A1(n_0_0_88), .A2(n_0_0_80), .ZN(n_23));
   NOR2_X1 i_0_0_145 (.A1(n_0_0_9), .A2(1'b0), .ZN(n_0_0_89));
   NAND2_X1 i_0_0_146 (.A1(n_0_0_73), .A2(n_0_0_89), .ZN(n_0_0_90));
   NOR2_X1 i_0_0_147 (.A1(n_0_0_71), .A2(n_0_0_90), .ZN(n_24));
   NAND2_X1 i_0_0_148 (.A1(n_0_0_76), .A2(n_0_0_89), .ZN(n_0_0_91));
   NOR2_X1 i_0_0_149 (.A1(n_0_0_71), .A2(n_0_0_91), .ZN(n_25));
   NAND2_X1 i_0_0_150 (.A1(n_0_0_78), .A2(n_0_0_89), .ZN(n_0_0_92));
   NOR2_X1 i_0_0_151 (.A1(n_0_0_71), .A2(n_0_0_92), .ZN(n_26));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_89), .A2(n_0_0_13), .ZN(n_0_0_93));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_71), .A2(n_0_0_93), .ZN(n_27));
   NOR2_X1 i_0_0_154 (.A1(n_0_0_81), .A2(n_0_0_90), .ZN(n_28));
   NOR2_X1 i_0_0_155 (.A1(n_0_0_81), .A2(n_0_0_91), .ZN(n_29));
   NOR2_X1 i_0_0_156 (.A1(n_0_0_81), .A2(n_0_0_92), .ZN(n_30));
   NOR2_X1 i_0_0_157 (.A1(n_0_0_81), .A2(n_0_0_93), .ZN(n_31));
   NOR2_X1 i_0_0_158 (.A1(1'b0), .A2(1'b0), .ZN(n_0_0_94));
   NAND2_X1 i_0_0_159 (.A1(n_0_0_73), .A2(n_0_0_94), .ZN(n_0_0_95));
   NOR2_X1 i_0_0_160 (.A1(n_0_0_71), .A2(n_0_0_95), .ZN(n_32));
   NAND2_X1 i_0_0_161 (.A1(n_0_0_76), .A2(n_0_0_94), .ZN(n_0_0_96));
   NOR2_X1 i_0_0_162 (.A1(n_0_0_71), .A2(n_0_0_96), .ZN(n_33));
   NAND2_X1 i_0_0_163 (.A1(n_0_0_78), .A2(n_0_0_94), .ZN(n_0_0_97));
   NOR2_X1 i_0_0_164 (.A1(n_0_0_71), .A2(n_0_0_97), .ZN(n_34));
   NAND2_X1 i_0_0_165 (.A1(n_0_0_13), .A2(n_0_0_94), .ZN(n_0_0_98));
   NOR2_X1 i_0_0_166 (.A1(n_0_0_71), .A2(n_0_0_98), .ZN(n_35));
   NOR2_X1 i_0_0_167 (.A1(n_0_0_81), .A2(n_0_0_95), .ZN(n_36));
   NOR2_X1 i_0_0_168 (.A1(n_0_0_81), .A2(n_0_0_96), .ZN(n_37));
   NOR2_X1 i_0_0_169 (.A1(n_0_0_81), .A2(n_0_0_97), .ZN(n_38));
   NOR2_X1 i_0_0_170 (.A1(n_0_0_81), .A2(n_0_0_98), .ZN(n_39));
   NOR2_X1 i_0_0_171 (.A1(n_0_0_82), .A2(n_0_0_90), .ZN(n_40));
   NOR2_X1 i_0_0_172 (.A1(n_0_0_82), .A2(n_0_0_91), .ZN(n_41));
   NOR2_X1 i_0_0_173 (.A1(n_0_0_82), .A2(n_0_0_92), .ZN(n_42));
   NOR2_X1 i_0_0_174 (.A1(n_0_0_82), .A2(n_0_0_93), .ZN(n_43));
   NOR2_X1 i_0_0_175 (.A1(n_0_0_88), .A2(n_0_0_90), .ZN(n_44));
   NOR2_X1 i_0_0_176 (.A1(n_0_0_88), .A2(n_0_0_91), .ZN(n_45));
   NOR2_X1 i_0_0_177 (.A1(n_0_0_88), .A2(n_0_0_92), .ZN(n_46));
   NOR2_X1 i_0_0_178 (.A1(n_0_0_88), .A2(n_0_0_93), .ZN(n_47));
   NOR2_X1 i_0_0_179 (.A1(n_0_0_82), .A2(n_0_0_95), .ZN(n_48));
   NOR2_X1 i_0_0_180 (.A1(n_0_0_82), .A2(n_0_0_96), .ZN(n_49));
   NOR2_X1 i_0_0_181 (.A1(n_0_0_82), .A2(n_0_0_97), .ZN(n_50));
   NOR2_X1 i_0_0_182 (.A1(n_0_0_82), .A2(n_0_0_98), .ZN(n_51));
   NOR2_X1 i_0_0_183 (.A1(n_0_0_88), .A2(n_0_0_95), .ZN(n_52));
   NOR2_X1 i_0_0_184 (.A1(n_0_0_88), .A2(n_0_0_96), .ZN(n_53));
   NOR2_X1 i_0_0_185 (.A1(n_0_0_88), .A2(n_0_0_97), .ZN(n_54));
   NOR2_X1 i_0_0_186 (.A1(n_0_0_88), .A2(n_0_0_98), .ZN(n_55));
   NOR2_X1 i_0_0_187 (.A1(n_0_0_69), .A2(1'b0), .ZN(n_0_0_99));
   NAND3_X1 i_0_0_188 (.A1(n_0_0_99), .A2(1'b0), .A3(1'b0), .ZN(n_0_0_100));
   NOR2_X1 i_0_0_189 (.A1(n_0_0_100), .A2(n_0_0_84), .ZN(n_56));
   NOR2_X1 i_0_0_190 (.A1(n_0_0_100), .A2(n_0_0_85), .ZN(n_57));
   NOR2_X1 i_0_0_191 (.A1(n_0_0_100), .A2(n_0_0_86), .ZN(n_58));
   NOR2_X1 i_0_0_192 (.A1(n_0_0_100), .A2(n_0_0_87), .ZN(n_59));
   NAND3_X1 i_0_0_193 (.A1(n_0_0_99), .A2(1'b0), .A3(n_0_0_8), .ZN(n_0_0_101));
   NOR2_X1 i_0_0_194 (.A1(n_0_0_101), .A2(n_0_0_84), .ZN(n_60));
   NOR2_X1 i_0_0_195 (.A1(n_0_0_101), .A2(n_0_0_85), .ZN(n_61));
   NOR2_X1 i_0_0_196 (.A1(n_0_0_101), .A2(n_0_0_86), .ZN(n_62));
   NOR2_X1 i_0_0_197 (.A1(n_0_0_101), .A2(n_0_0_87), .ZN(n_63));
   NOR2_X1 i_0_0_198 (.A1(n_0_0_100), .A2(n_0_0_75), .ZN(n_64));
   NOR2_X1 i_0_0_199 (.A1(n_0_0_100), .A2(n_0_0_77), .ZN(n_65));
   NOR2_X1 i_0_0_200 (.A1(n_0_0_100), .A2(n_0_0_79), .ZN(n_66));
   NOR2_X1 i_0_0_201 (.A1(n_0_0_100), .A2(n_0_0_80), .ZN(n_67));
   NOR2_X1 i_0_0_202 (.A1(n_0_0_101), .A2(n_0_0_75), .ZN(n_68));
   NOR2_X1 i_0_0_203 (.A1(n_0_0_101), .A2(n_0_0_77), .ZN(n_69));
   NOR2_X1 i_0_0_204 (.A1(n_0_0_101), .A2(n_0_0_79), .ZN(n_70));
   NOR2_X1 i_0_0_205 (.A1(n_0_0_101), .A2(n_0_0_80), .ZN(n_71));
   NAND3_X1 i_0_0_206 (.A1(n_0_0_99), .A2(n_0_0_3), .A3(1'b0), .ZN(n_0_0_102));
   NOR2_X1 i_0_0_207 (.A1(n_0_0_102), .A2(n_0_0_84), .ZN(n_72));
   NOR2_X1 i_0_0_208 (.A1(n_0_0_102), .A2(n_0_0_85), .ZN(n_73));
   NOR2_X1 i_0_0_209 (.A1(n_0_0_102), .A2(n_0_0_86), .ZN(n_74));
   NOR2_X1 i_0_0_210 (.A1(n_0_0_102), .A2(n_0_0_87), .ZN(n_75));
   NAND3_X1 i_0_0_211 (.A1(n_0_0_99), .A2(n_0_0_3), .A3(n_0_0_8), .ZN(n_0_0_103));
   NOR2_X1 i_0_0_212 (.A1(n_0_0_103), .A2(n_0_0_84), .ZN(n_76));
   NOR2_X1 i_0_0_213 (.A1(n_0_0_103), .A2(n_0_0_85), .ZN(n_77));
   NOR2_X1 i_0_0_214 (.A1(n_0_0_103), .A2(n_0_0_86), .ZN(n_78));
   NOR2_X1 i_0_0_215 (.A1(n_0_0_103), .A2(n_0_0_87), .ZN(n_79));
   NOR2_X1 i_0_0_216 (.A1(n_0_0_102), .A2(n_0_0_75), .ZN(n_80));
   NOR2_X1 i_0_0_217 (.A1(n_0_0_102), .A2(n_0_0_77), .ZN(n_81));
   NOR2_X1 i_0_0_218 (.A1(n_0_0_102), .A2(n_0_0_79), .ZN(n_82));
   NOR2_X1 i_0_0_219 (.A1(n_0_0_102), .A2(n_0_0_80), .ZN(n_83));
   NOR2_X1 i_0_0_220 (.A1(n_0_0_103), .A2(n_0_0_75), .ZN(n_84));
   NOR2_X1 i_0_0_221 (.A1(n_0_0_103), .A2(n_0_0_77), .ZN(n_85));
   NOR2_X1 i_0_0_222 (.A1(n_0_0_103), .A2(n_0_0_79), .ZN(n_86));
   NOR2_X1 i_0_0_223 (.A1(n_0_0_103), .A2(n_0_0_80), .ZN(n_87));
   NOR2_X1 i_0_0_224 (.A1(n_0_0_100), .A2(n_0_0_90), .ZN(n_88));
   NOR2_X1 i_0_0_225 (.A1(n_0_0_100), .A2(n_0_0_91), .ZN(n_89));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_100), .A2(n_0_0_92), .ZN(n_90));
   NOR2_X1 i_0_0_227 (.A1(n_0_0_100), .A2(n_0_0_93), .ZN(n_91));
   NOR2_X1 i_0_0_228 (.A1(n_0_0_101), .A2(n_0_0_90), .ZN(n_92));
   NOR2_X1 i_0_0_229 (.A1(n_0_0_101), .A2(n_0_0_91), .ZN(n_93));
   NOR2_X1 i_0_0_230 (.A1(n_0_0_101), .A2(n_0_0_92), .ZN(n_94));
   NOR2_X1 i_0_0_231 (.A1(n_0_0_101), .A2(n_0_0_93), .ZN(n_95));
   NOR2_X1 i_0_0_232 (.A1(n_0_0_100), .A2(n_0_0_95), .ZN(n_96));
   NOR2_X1 i_0_0_233 (.A1(n_0_0_100), .A2(n_0_0_96), .ZN(n_97));
   NOR2_X1 i_0_0_234 (.A1(n_0_0_100), .A2(n_0_0_97), .ZN(n_98));
   NOR2_X1 i_0_0_235 (.A1(n_0_0_100), .A2(n_0_0_98), .ZN(n_99));
   NOR2_X1 i_0_0_236 (.A1(n_0_0_101), .A2(n_0_0_95), .ZN(n_100));
   NOR2_X1 i_0_0_237 (.A1(n_0_0_101), .A2(n_0_0_96), .ZN(n_101));
   NOR2_X1 i_0_0_238 (.A1(n_0_0_101), .A2(n_0_0_97), .ZN(n_102));
   NOR2_X1 i_0_0_239 (.A1(n_0_0_101), .A2(n_0_0_98), .ZN(n_103));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_102), .A2(n_0_0_90), .ZN(n_104));
   NOR2_X1 i_0_0_241 (.A1(n_0_0_102), .A2(n_0_0_91), .ZN(n_105));
   NOR2_X1 i_0_0_242 (.A1(n_0_0_102), .A2(n_0_0_92), .ZN(n_106));
   NOR2_X1 i_0_0_243 (.A1(n_0_0_102), .A2(n_0_0_93), .ZN(n_107));
   NOR2_X1 i_0_0_244 (.A1(n_0_0_103), .A2(n_0_0_90), .ZN(n_108));
   NOR2_X1 i_0_0_245 (.A1(n_0_0_103), .A2(n_0_0_91), .ZN(n_109));
   NOR2_X1 i_0_0_246 (.A1(n_0_0_103), .A2(n_0_0_92), .ZN(n_110));
   NOR2_X1 i_0_0_247 (.A1(n_0_0_103), .A2(n_0_0_93), .ZN(n_111));
   NOR2_X1 i_0_0_248 (.A1(n_0_0_102), .A2(n_0_0_95), .ZN(n_112));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_102), .A2(n_0_0_96), .ZN(n_113));
   NOR2_X1 i_0_0_250 (.A1(n_0_0_102), .A2(n_0_0_97), .ZN(n_114));
   NOR2_X1 i_0_0_251 (.A1(n_0_0_102), .A2(n_0_0_98), .ZN(n_115));
   NOR2_X1 i_0_0_252 (.A1(n_0_0_103), .A2(n_0_0_95), .ZN(n_116));
   NOR2_X1 i_0_0_253 (.A1(n_0_0_103), .A2(n_0_0_96), .ZN(n_117));
   NOR2_X1 i_0_0_254 (.A1(n_0_0_103), .A2(n_0_0_97), .ZN(n_118));
   NOR2_X1 i_0_0_255 (.A1(n_0_0_103), .A2(n_0_0_98), .ZN(n_119));
   INV_X1 i_0_0_256 (.A(clk), .ZN(n_120));
   DFF_X1 \address_reg[9]  (.D(i_address[9]), .CK(n_1_0), .Q(o_mem_addr[9]), 
      .QN());
   DFF_X1 \address_reg[8]  (.D(i_address[8]), .CK(n_1_0), .Q(o_mem_addr[8]), 
      .QN());
   DFF_X1 \address_reg[7]  (.D(i_address[7]), .CK(n_1_0), .Q(o_mem_addr[7]), 
      .QN());
   DFF_X1 \address_reg[6]  (.D(i_address[6]), .CK(n_1_0), .Q(o_mem_addr[6]), 
      .QN());
   DFF_X1 \address_reg[5]  (.D(i_address[5]), .CK(n_1_0), .Q(o_mem_addr[5]), 
      .QN());
   DFF_X1 \address_reg[4]  (.D(i_address[4]), .CK(n_1_0), .Q(o_mem_addr[4]), 
      .QN());
   DFF_X1 \address_reg[3]  (.D(i_address[3]), .CK(n_1_0), .Q(o_mem_addr[3]), 
      .QN());
   DFF_X1 \address_reg[2]  (.D(i_address[2]), .CK(n_1_0), .Q(o_mem_addr[2]), 
      .QN());
   DFF_X1 \address_reg[1]  (.D(i_address[1]), .CK(n_1_0), .Q(o_mem_addr[1]), 
      .QN());
   DFF_X1 \address_reg[0]  (.D(i_address[0]), .CK(n_1_0), .Q(o_mem_addr[0]), 
      .QN());
   DFF_X1 read_reg (.D(n_1_3), .CK(clk), .Q(read), .QN());
   MUX2_X1 read_reg_enable_mux_0 (.A(read), .B(n_1_2), .S(n_1_1), .Z(n_1_3));
   DFF_X1 \count_reg[9]  (.D(i_count[9]), .CK(n_1_0), .Q(count[9]), .QN());
   DFF_X1 \count_reg[8]  (.D(i_count[8]), .CK(n_1_0), .Q(count[8]), .QN());
   DFF_X1 \count_reg[7]  (.D(i_count[7]), .CK(n_1_0), .Q(count[7]), .QN());
   DFF_X1 \count_reg[6]  (.D(i_count[6]), .CK(n_1_0), .Q(count[6]), .QN());
   DFF_X1 \count_reg[5]  (.D(i_count[5]), .CK(n_1_0), .Q(count[5]), .QN());
   DFF_X1 \count_reg[4]  (.D(i_count[4]), .CK(n_1_0), .Q(count[4]), .QN());
   DFF_X1 \count_reg[3]  (.D(i_count[3]), .CK(n_1_0), .Q(count[3]), .QN());
   DFF_X1 \count_reg[2]  (.D(i_count[2]), .CK(n_1_0), .Q(count[2]), .QN());
   DFF_X1 \count_reg[1]  (.D(i_count[1]), .CK(n_1_0), .Q(count[1]), .QN());
   DFF_X1 \count_reg[0]  (.D(i_count[0]), .CK(n_1_0), .Q(count[0]), .QN());
   CLKGATETST_X1 clk_gate_count_reg (.CK(clk), .E(n_1_2), .SE(1'b0), .GCK(n_1_0));
   OAI21_X1 i_1_0_0 (.A(n_1_0_0), .B1(n_1_0_4), .B2(read), .ZN(n_1_1));
   NAND4_X1 i_1_0_1 (.A1(read), .A2(n_1_0_3), .A3(n_1_0_2), .A4(n_1_0_1), 
      .ZN(n_1_0_0));
   NOR4_X1 i_1_0_2 (.A1(count[8]), .A2(count[7]), .A3(count[5]), .A4(count[2]), 
      .ZN(n_1_0_1));
   NOR4_X1 i_1_0_3 (.A1(count[9]), .A2(count[6]), .A3(count[4]), .A4(count[3]), 
      .ZN(n_1_0_2));
   NOR2_X1 i_1_0_4 (.A1(count[1]), .A2(count[0]), .ZN(n_1_0_3));
   NOR2_X1 i_1_0_5 (.A1(n_1_0_4), .A2(read), .ZN(n_1_2));
   INV_X1 i_1_0_6 (.A(i_read), .ZN(n_1_0_4));
endmodule
