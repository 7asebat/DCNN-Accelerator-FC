/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 04:51:33 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3896383824 */

module Softmax(\values[0] , \values[1] , \values[2] , \values[3] , \values[4] , 
      \values[5] , \values[6] , \values[7] , \values[8] , \values[9] , class_out);
   input [15:0]\values[0] ;
   input [15:0]\values[1] ;
   input [15:0]\values[2] ;
   input [15:0]\values[3] ;
   input [15:0]\values[4] ;
   input [15:0]\values[5] ;
   input [15:0]\values[6] ;
   input [15:0]\values[7] ;
   input [15:0]\values[8] ;
   input [15:0]\values[9] ;
   output [15:0]class_out;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;

   assign class_out[15] = class_out[4];
   assign class_out[14] = class_out[4];
   assign class_out[13] = class_out[4];
   assign class_out[12] = class_out[4];
   assign class_out[11] = class_out[4];
   assign class_out[10] = class_out[4];
   assign class_out[9] = class_out[4];
   assign class_out[8] = class_out[4];
   assign class_out[7] = class_out[4];
   assign class_out[6] = class_out[4];
   assign class_out[5] = class_out[4];

   NAND2_X1 i_0_0_0 (.A1(n_0_0_8), .A2(n_0_0_0), .ZN(class_out[0]));
   OAI21_X1 i_0_0_1 (.A(n_0_0_64), .B1(n_0_0_1), .B2(n_0_0_121), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_2), .ZN(n_0_0_1));
   OAI21_X1 i_0_0_3 (.A(n_0_0_178), .B1(n_0_0_3), .B2(n_0_0_238), .ZN(n_0_0_2));
   AOI21_X1 i_0_0_4 (.A(n_0_0_292), .B1(n_0_0_4), .B2(n_0_0_355), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_5 (.A(n_0_0_417), .B1(n_0_0_349), .B2(n_0_0_479), .ZN(n_0_0_4));
   AOI21_X1 i_0_0_6 (.A(n_0_0_6), .B1(n_0_0_5), .B2(n_0_0_120), .ZN(class_out[1]));
   OAI21_X1 i_0_0_7 (.A(n_0_0_237), .B1(n_0_0_347), .B2(n_0_0_354), .ZN(n_0_0_5));
   AOI21_X1 i_0_0_8 (.A(n_0_0_6), .B1(n_0_0_119), .B2(n_0_0_345), .ZN(
      class_out[2]));
   NAND2_X1 i_0_0_9 (.A1(n_0_0_7), .A2(n_0_0_118), .ZN(class_out[3]));
   NOR2_X1 i_0_0_10 (.A1(n_0_0_118), .A2(n_0_0_6), .ZN(class_out[4]));
   INV_X1 i_0_0_11 (.A(n_0_0_7), .ZN(n_0_0_6));
   AOI21_X1 i_0_0_12 (.A(n_0_0_9), .B1(n_0_0_65), .B2(n_0_0_66), .ZN(n_0_0_7));
   INV_X1 i_0_0_13 (.A(n_0_0_9), .ZN(n_0_0_8));
   AOI22_X1 i_0_0_14 (.A1(n_0_0_12), .A2(n_0_0_10), .B1(\values[9] [15]), 
      .B2(n_0_0_63), .ZN(n_0_0_9));
   AOI21_X1 i_0_0_15 (.A(n_0_0_11), .B1(n_0_0_13), .B2(\values[9] [14]), 
      .ZN(n_0_0_10));
   NOR2_X1 i_0_0_16 (.A1(n_0_0_63), .A2(\values[9] [15]), .ZN(n_0_0_11));
   OAI21_X1 i_0_0_17 (.A(n_0_0_15), .B1(n_0_0_13), .B2(\values[9] [14]), 
      .ZN(n_0_0_12));
   OAI21_X1 i_0_0_18 (.A(n_0_0_14), .B1(n_0_0_64), .B2(\values[8] [14]), 
      .ZN(n_0_0_13));
   NAND2_X1 i_0_0_19 (.A1(n_0_0_70), .A2(n_0_0_64), .ZN(n_0_0_14));
   OAI21_X1 i_0_0_20 (.A(n_0_0_16), .B1(n_0_0_20), .B2(n_0_0_17), .ZN(n_0_0_15));
   NAND2_X1 i_0_0_21 (.A1(\values[9] [13]), .A2(n_0_0_18), .ZN(n_0_0_16));
   OAI22_X1 i_0_0_22 (.A1(\values[9] [12]), .A2(n_0_0_21), .B1(n_0_0_18), 
      .B2(\values[9] [13]), .ZN(n_0_0_17));
   OAI21_X1 i_0_0_23 (.A(n_0_0_19), .B1(n_0_0_64), .B2(\values[8] [13]), 
      .ZN(n_0_0_18));
   NAND2_X1 i_0_0_24 (.A1(n_0_0_74), .A2(n_0_0_64), .ZN(n_0_0_19));
   AOI221_X1 i_0_0_25 (.A(n_0_0_23), .B1(n_0_0_21), .B2(\values[9] [12]), 
      .C1(\values[9] [11]), .C2(n_0_0_25), .ZN(n_0_0_20));
   OAI21_X1 i_0_0_26 (.A(n_0_0_22), .B1(n_0_0_64), .B2(\values[8] [12]), 
      .ZN(n_0_0_21));
   NAND2_X1 i_0_0_27 (.A1(n_0_0_77), .A2(n_0_0_64), .ZN(n_0_0_22));
   AOI21_X1 i_0_0_28 (.A(n_0_0_24), .B1(n_0_0_30), .B2(n_0_0_27), .ZN(n_0_0_23));
   OAI22_X1 i_0_0_29 (.A1(\values[9] [10]), .A2(n_0_0_28), .B1(n_0_0_25), 
      .B2(\values[9] [11]), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_30 (.A(n_0_0_26), .B1(n_0_0_64), .B2(\values[8] [11]), 
      .ZN(n_0_0_25));
   NAND2_X1 i_0_0_31 (.A1(n_0_0_80), .A2(n_0_0_64), .ZN(n_0_0_26));
   AOI22_X1 i_0_0_32 (.A1(\values[9] [9]), .A2(n_0_0_31), .B1(n_0_0_28), 
      .B2(\values[9] [10]), .ZN(n_0_0_27));
   OAI21_X1 i_0_0_33 (.A(n_0_0_29), .B1(n_0_0_64), .B2(\values[8] [10]), 
      .ZN(n_0_0_28));
   NAND2_X1 i_0_0_34 (.A1(n_0_0_84), .A2(n_0_0_64), .ZN(n_0_0_29));
   OAI221_X1 i_0_0_35 (.A(n_0_0_33), .B1(n_0_0_31), .B2(\values[9] [9]), 
      .C1(\values[9] [8]), .C2(n_0_0_35), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_36 (.A(n_0_0_32), .B1(n_0_0_64), .B2(\values[8] [9]), .ZN(
      n_0_0_31));
   NAND2_X1 i_0_0_37 (.A1(n_0_0_87), .A2(n_0_0_64), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_38 (.A(n_0_0_34), .B1(n_0_0_40), .B2(n_0_0_37), .ZN(n_0_0_33));
   AOI22_X1 i_0_0_39 (.A1(\values[9] [7]), .A2(n_0_0_38), .B1(n_0_0_35), 
      .B2(\values[9] [8]), .ZN(n_0_0_34));
   OAI21_X1 i_0_0_40 (.A(n_0_0_36), .B1(n_0_0_64), .B2(\values[8] [8]), .ZN(
      n_0_0_35));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_90), .A2(n_0_0_64), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_42 (.A1(\values[9] [6]), .A2(n_0_0_41), .B1(n_0_0_38), 
      .B2(\values[9] [7]), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_43 (.A(n_0_0_39), .B1(n_0_0_64), .B2(\values[8] [7]), .ZN(
      n_0_0_38));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_94), .A2(n_0_0_64), .ZN(n_0_0_39));
   AOI221_X1 i_0_0_45 (.A(n_0_0_44), .B1(n_0_0_41), .B2(\values[9] [6]), 
      .C1(\values[9] [5]), .C2(n_0_0_46), .ZN(n_0_0_40));
   INV_X1 i_0_0_46 (.A(n_0_0_42), .ZN(n_0_0_41));
   AOI21_X1 i_0_0_47 (.A(n_0_0_43), .B1(n_0_0_64), .B2(n_0_0_97), .ZN(n_0_0_42));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_64), .A2(\values[8] [6]), .ZN(n_0_0_43));
   AOI21_X1 i_0_0_49 (.A(n_0_0_45), .B1(n_0_0_51), .B2(n_0_0_48), .ZN(n_0_0_44));
   OAI22_X1 i_0_0_50 (.A1(\values[9] [4]), .A2(n_0_0_49), .B1(n_0_0_46), 
      .B2(\values[9] [5]), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_51 (.A(n_0_0_47), .B1(n_0_0_64), .B2(\values[8] [5]), .ZN(
      n_0_0_46));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_100), .A2(n_0_0_64), .ZN(n_0_0_47));
   AOI22_X1 i_0_0_53 (.A1(\values[9] [3]), .A2(n_0_0_52), .B1(n_0_0_49), 
      .B2(\values[9] [4]), .ZN(n_0_0_48));
   OAI21_X1 i_0_0_54 (.A(n_0_0_50), .B1(n_0_0_64), .B2(\values[8] [4]), .ZN(
      n_0_0_49));
   NAND2_X1 i_0_0_55 (.A1(n_0_0_104), .A2(n_0_0_64), .ZN(n_0_0_50));
   OAI221_X1 i_0_0_56 (.A(n_0_0_54), .B1(n_0_0_52), .B2(\values[9] [3]), 
      .C1(\values[9] [2]), .C2(n_0_0_56), .ZN(n_0_0_51));
   OAI21_X1 i_0_0_57 (.A(n_0_0_53), .B1(n_0_0_64), .B2(\values[8] [3]), .ZN(
      n_0_0_52));
   NAND2_X1 i_0_0_58 (.A1(n_0_0_107), .A2(n_0_0_64), .ZN(n_0_0_53));
   OAI21_X1 i_0_0_59 (.A(n_0_0_55), .B1(n_0_0_58), .B2(n_0_0_59), .ZN(n_0_0_54));
   AOI22_X1 i_0_0_60 (.A1(\values[9] [1]), .A2(n_0_0_60), .B1(n_0_0_56), 
      .B2(\values[9] [2]), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_61 (.A(n_0_0_57), .B1(n_0_0_64), .B2(\values[8] [2]), .ZN(
      n_0_0_56));
   NAND2_X1 i_0_0_62 (.A1(n_0_0_111), .A2(n_0_0_64), .ZN(n_0_0_57));
   OAI221_X1 i_0_0_63 (.A(\values[9] [0]), .B1(n_0_0_64), .B2(n_0_0_506), 
      .C1(n_0_0_60), .C2(\values[9] [1]), .ZN(n_0_0_58));
   AND2_X1 i_0_0_64 (.A1(n_0_0_114), .A2(n_0_0_64), .ZN(n_0_0_59));
   INV_X1 i_0_0_65 (.A(n_0_0_61), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_66 (.A(n_0_0_62), .B1(n_0_0_64), .B2(n_0_0_507), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_67 (.A1(n_0_0_64), .A2(n_0_0_116), .ZN(n_0_0_62));
   NAND3_X1 i_0_0_68 (.A1(\values[7] [15]), .A2(\values[8] [15]), .A3(n_0_0_176), 
      .ZN(n_0_0_63));
   NAND2_X1 i_0_0_69 (.A1(n_0_0_66), .A2(n_0_0_65), .ZN(n_0_0_64));
   NAND2_X1 i_0_0_70 (.A1(n_0_0_68), .A2(\values[8] [15]), .ZN(n_0_0_65));
   OAI211_X1 i_0_0_71 (.A(n_0_0_69), .B(n_0_0_67), .C1(n_0_0_68), .C2(
      \values[8] [15]), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_72 (.A1(n_0_0_70), .A2(\values[8] [14]), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_73 (.A1(\values[7] [15]), .A2(n_0_0_176), .ZN(n_0_0_68));
   OAI221_X1 i_0_0_74 (.A(n_0_0_72), .B1(n_0_0_70), .B2(\values[8] [14]), 
      .C1(\values[8] [13]), .C2(n_0_0_74), .ZN(n_0_0_69));
   AOI21_X1 i_0_0_75 (.A(n_0_0_71), .B1(n_0_0_121), .B2(\values[7] [14]), 
      .ZN(n_0_0_70));
   NOR2_X1 i_0_0_76 (.A1(n_0_0_121), .A2(n_0_0_125), .ZN(n_0_0_71));
   OAI21_X1 i_0_0_77 (.A(n_0_0_73), .B1(n_0_0_79), .B2(n_0_0_76), .ZN(n_0_0_72));
   AOI22_X1 i_0_0_78 (.A1(\values[8] [12]), .A2(n_0_0_77), .B1(n_0_0_74), 
      .B2(\values[8] [13]), .ZN(n_0_0_73));
   AOI21_X1 i_0_0_79 (.A(n_0_0_75), .B1(n_0_0_121), .B2(\values[7] [13]), 
      .ZN(n_0_0_74));
   NOR2_X1 i_0_0_80 (.A1(n_0_0_121), .A2(n_0_0_129), .ZN(n_0_0_75));
   OAI22_X1 i_0_0_81 (.A1(\values[8] [11]), .A2(n_0_0_80), .B1(n_0_0_77), 
      .B2(\values[8] [12]), .ZN(n_0_0_76));
   AOI21_X1 i_0_0_82 (.A(n_0_0_78), .B1(n_0_0_121), .B2(\values[7] [12]), 
      .ZN(n_0_0_77));
   NOR2_X1 i_0_0_83 (.A1(n_0_0_121), .A2(n_0_0_132), .ZN(n_0_0_78));
   AOI221_X1 i_0_0_84 (.A(n_0_0_82), .B1(n_0_0_80), .B2(\values[8] [11]), 
      .C1(\values[8] [10]), .C2(n_0_0_84), .ZN(n_0_0_79));
   AOI21_X1 i_0_0_85 (.A(n_0_0_81), .B1(n_0_0_121), .B2(\values[7] [11]), 
      .ZN(n_0_0_80));
   NOR2_X1 i_0_0_86 (.A1(n_0_0_121), .A2(n_0_0_135), .ZN(n_0_0_81));
   AOI21_X1 i_0_0_87 (.A(n_0_0_83), .B1(n_0_0_89), .B2(n_0_0_86), .ZN(n_0_0_82));
   OAI22_X1 i_0_0_88 (.A1(\values[8] [9]), .A2(n_0_0_87), .B1(n_0_0_84), 
      .B2(\values[8] [10]), .ZN(n_0_0_83));
   AOI21_X1 i_0_0_89 (.A(n_0_0_85), .B1(n_0_0_121), .B2(\values[7] [10]), 
      .ZN(n_0_0_84));
   NOR2_X1 i_0_0_90 (.A1(n_0_0_121), .A2(n_0_0_139), .ZN(n_0_0_85));
   AOI22_X1 i_0_0_91 (.A1(\values[8] [8]), .A2(n_0_0_90), .B1(n_0_0_87), 
      .B2(\values[8] [9]), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_92 (.A(n_0_0_88), .B1(n_0_0_121), .B2(\values[7] [9]), 
      .ZN(n_0_0_87));
   NOR2_X1 i_0_0_93 (.A1(n_0_0_121), .A2(n_0_0_142), .ZN(n_0_0_88));
   OAI221_X1 i_0_0_94 (.A(n_0_0_92), .B1(n_0_0_90), .B2(\values[8] [8]), 
      .C1(\values[8] [7]), .C2(n_0_0_94), .ZN(n_0_0_89));
   AOI21_X1 i_0_0_95 (.A(n_0_0_91), .B1(n_0_0_121), .B2(\values[7] [8]), 
      .ZN(n_0_0_90));
   NOR2_X1 i_0_0_96 (.A1(n_0_0_121), .A2(n_0_0_173), .ZN(n_0_0_91));
   OAI21_X1 i_0_0_97 (.A(n_0_0_93), .B1(n_0_0_99), .B2(n_0_0_96), .ZN(n_0_0_92));
   AOI22_X1 i_0_0_98 (.A1(\values[8] [6]), .A2(n_0_0_97), .B1(n_0_0_94), 
      .B2(\values[8] [7]), .ZN(n_0_0_93));
   AOI21_X1 i_0_0_99 (.A(n_0_0_95), .B1(n_0_0_121), .B2(\values[7] [7]), 
      .ZN(n_0_0_94));
   NOR2_X1 i_0_0_100 (.A1(n_0_0_121), .A2(n_0_0_148), .ZN(n_0_0_95));
   OAI22_X1 i_0_0_101 (.A1(\values[8] [5]), .A2(n_0_0_100), .B1(n_0_0_97), 
      .B2(\values[8] [6]), .ZN(n_0_0_96));
   AOI21_X1 i_0_0_102 (.A(n_0_0_98), .B1(n_0_0_121), .B2(\values[7] [6]), 
      .ZN(n_0_0_97));
   NOR2_X1 i_0_0_103 (.A1(n_0_0_121), .A2(n_0_0_151), .ZN(n_0_0_98));
   AOI221_X1 i_0_0_104 (.A(n_0_0_102), .B1(n_0_0_100), .B2(\values[8] [5]), 
      .C1(\values[8] [4]), .C2(n_0_0_104), .ZN(n_0_0_99));
   AOI21_X1 i_0_0_105 (.A(n_0_0_101), .B1(n_0_0_121), .B2(\values[7] [5]), 
      .ZN(n_0_0_100));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_121), .A2(n_0_0_155), .ZN(n_0_0_101));
   AOI21_X1 i_0_0_107 (.A(n_0_0_103), .B1(n_0_0_109), .B2(n_0_0_106), .ZN(
      n_0_0_102));
   OAI22_X1 i_0_0_108 (.A1(\values[8] [3]), .A2(n_0_0_107), .B1(n_0_0_104), 
      .B2(\values[8] [4]), .ZN(n_0_0_103));
   AOI21_X1 i_0_0_109 (.A(n_0_0_105), .B1(n_0_0_121), .B2(\values[7] [4]), 
      .ZN(n_0_0_104));
   NOR2_X1 i_0_0_110 (.A1(n_0_0_121), .A2(n_0_0_158), .ZN(n_0_0_105));
   AOI22_X1 i_0_0_111 (.A1(\values[8] [2]), .A2(n_0_0_111), .B1(n_0_0_107), 
      .B2(\values[8] [3]), .ZN(n_0_0_106));
   AOI21_X1 i_0_0_112 (.A(n_0_0_108), .B1(n_0_0_121), .B2(\values[7] [3]), 
      .ZN(n_0_0_107));
   NOR2_X1 i_0_0_113 (.A1(n_0_0_121), .A2(n_0_0_171), .ZN(n_0_0_108));
   OAI211_X1 i_0_0_114 (.A(n_0_0_113), .B(n_0_0_110), .C1(n_0_0_111), .C2(
      \values[8] [2]), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_115 (.A1(n_0_0_116), .A2(n_0_0_507), .ZN(n_0_0_110));
   AOI21_X1 i_0_0_116 (.A(n_0_0_112), .B1(n_0_0_121), .B2(\values[7] [2]), 
      .ZN(n_0_0_111));
   NOR2_X1 i_0_0_117 (.A1(n_0_0_121), .A2(n_0_0_169), .ZN(n_0_0_112));
   OAI22_X1 i_0_0_118 (.A1(n_0_0_507), .A2(n_0_0_116), .B1(n_0_0_114), .B2(
      n_0_0_506), .ZN(n_0_0_113));
   OAI21_X1 i_0_0_119 (.A(n_0_0_115), .B1(n_0_0_121), .B2(n_0_0_166), .ZN(
      n_0_0_114));
   NAND2_X1 i_0_0_120 (.A1(n_0_0_121), .A2(\values[7] [0]), .ZN(n_0_0_115));
   OAI21_X1 i_0_0_121 (.A(n_0_0_117), .B1(n_0_0_121), .B2(n_0_0_164), .ZN(
      n_0_0_116));
   NAND2_X1 i_0_0_122 (.A1(n_0_0_121), .A2(\values[7] [1]), .ZN(n_0_0_117));
   NAND2_X1 i_0_0_123 (.A1(n_0_0_346), .A2(n_0_0_119), .ZN(n_0_0_118));
   AND2_X1 i_0_0_124 (.A1(n_0_0_237), .A2(n_0_0_120), .ZN(n_0_0_119));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_121), .A2(n_0_0_177), .ZN(n_0_0_120));
   OAI22_X1 i_0_0_126 (.A1(n_0_0_122), .A2(n_0_0_124), .B1(n_0_0_175), .B2(
      \values[7] [15]), .ZN(n_0_0_121));
   OAI21_X1 i_0_0_127 (.A(n_0_0_123), .B1(n_0_0_125), .B2(\values[7] [14]), 
      .ZN(n_0_0_122));
   NAND2_X1 i_0_0_128 (.A1(n_0_0_175), .A2(\values[7] [15]), .ZN(n_0_0_123));
   AOI221_X1 i_0_0_129 (.A(n_0_0_127), .B1(n_0_0_125), .B2(\values[7] [14]), 
      .C1(\values[7] [13]), .C2(n_0_0_129), .ZN(n_0_0_124));
   OAI21_X1 i_0_0_130 (.A(n_0_0_126), .B1(n_0_0_178), .B2(\values[6] [14]), 
      .ZN(n_0_0_125));
   NAND2_X1 i_0_0_131 (.A1(n_0_0_234), .A2(n_0_0_178), .ZN(n_0_0_126));
   AOI21_X1 i_0_0_132 (.A(n_0_0_128), .B1(n_0_0_134), .B2(n_0_0_131), .ZN(
      n_0_0_127));
   OAI22_X1 i_0_0_133 (.A1(\values[7] [12]), .A2(n_0_0_132), .B1(n_0_0_129), 
      .B2(\values[7] [13]), .ZN(n_0_0_128));
   OAI21_X1 i_0_0_134 (.A(n_0_0_130), .B1(n_0_0_178), .B2(\values[6] [13]), 
      .ZN(n_0_0_129));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_230), .A2(n_0_0_178), .ZN(n_0_0_130));
   AOI22_X1 i_0_0_136 (.A1(\values[7] [11]), .A2(n_0_0_135), .B1(n_0_0_132), 
      .B2(\values[7] [12]), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_137 (.A(n_0_0_133), .B1(n_0_0_178), .B2(\values[6] [12]), 
      .ZN(n_0_0_132));
   NAND2_X1 i_0_0_138 (.A1(n_0_0_228), .A2(n_0_0_178), .ZN(n_0_0_133));
   OAI221_X1 i_0_0_139 (.A(n_0_0_137), .B1(n_0_0_135), .B2(\values[7] [11]), 
      .C1(\values[7] [10]), .C2(n_0_0_139), .ZN(n_0_0_134));
   OAI21_X1 i_0_0_140 (.A(n_0_0_136), .B1(n_0_0_178), .B2(\values[6] [11]), 
      .ZN(n_0_0_135));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_190), .A2(n_0_0_178), .ZN(n_0_0_136));
   OAI21_X1 i_0_0_142 (.A(n_0_0_138), .B1(n_0_0_141), .B2(n_0_0_144), .ZN(
      n_0_0_137));
   AOI22_X1 i_0_0_143 (.A1(\values[7] [9]), .A2(n_0_0_142), .B1(n_0_0_139), 
      .B2(\values[7] [10]), .ZN(n_0_0_138));
   OAI21_X1 i_0_0_144 (.A(n_0_0_140), .B1(n_0_0_178), .B2(\values[6] [10]), 
      .ZN(n_0_0_139));
   NAND2_X1 i_0_0_145 (.A1(n_0_0_193), .A2(n_0_0_178), .ZN(n_0_0_140));
   NOR2_X1 i_0_0_146 (.A1(\values[7] [9]), .A2(n_0_0_142), .ZN(n_0_0_141));
   OAI21_X1 i_0_0_147 (.A(n_0_0_143), .B1(n_0_0_178), .B2(\values[6] [9]), 
      .ZN(n_0_0_142));
   NAND2_X1 i_0_0_148 (.A1(n_0_0_197), .A2(n_0_0_178), .ZN(n_0_0_143));
   AOI21_X1 i_0_0_149 (.A(n_0_0_145), .B1(n_0_0_173), .B2(\values[7] [8]), 
      .ZN(n_0_0_144));
   AOI21_X1 i_0_0_150 (.A(n_0_0_146), .B1(n_0_0_150), .B2(n_0_0_147), .ZN(
      n_0_0_145));
   OAI22_X1 i_0_0_151 (.A1(\values[7] [8]), .A2(n_0_0_173), .B1(n_0_0_148), 
      .B2(\values[7] [7]), .ZN(n_0_0_146));
   AOI22_X1 i_0_0_152 (.A1(\values[7] [6]), .A2(n_0_0_151), .B1(n_0_0_148), 
      .B2(\values[7] [7]), .ZN(n_0_0_147));
   OAI21_X1 i_0_0_153 (.A(n_0_0_149), .B1(n_0_0_178), .B2(\values[6] [7]), 
      .ZN(n_0_0_148));
   NAND2_X1 i_0_0_154 (.A1(n_0_0_178), .A2(n_0_0_203), .ZN(n_0_0_149));
   OAI221_X1 i_0_0_155 (.A(n_0_0_153), .B1(n_0_0_151), .B2(\values[7] [6]), 
      .C1(\values[7] [5]), .C2(n_0_0_155), .ZN(n_0_0_150));
   OAI21_X1 i_0_0_156 (.A(n_0_0_152), .B1(n_0_0_178), .B2(\values[6] [6]), 
      .ZN(n_0_0_151));
   NAND2_X1 i_0_0_157 (.A1(n_0_0_178), .A2(n_0_0_207), .ZN(n_0_0_152));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_157), .A2(n_0_0_154), .ZN(n_0_0_153));
   AOI22_X1 i_0_0_159 (.A1(\values[7] [4]), .A2(n_0_0_158), .B1(n_0_0_155), 
      .B2(\values[7] [5]), .ZN(n_0_0_154));
   OAI21_X1 i_0_0_160 (.A(n_0_0_156), .B1(n_0_0_178), .B2(\values[6] [5]), 
      .ZN(n_0_0_155));
   NAND2_X1 i_0_0_161 (.A1(n_0_0_178), .A2(n_0_0_210), .ZN(n_0_0_156));
   OAI221_X1 i_0_0_162 (.A(n_0_0_160), .B1(n_0_0_158), .B2(\values[7] [4]), 
      .C1(\values[7] [3]), .C2(n_0_0_171), .ZN(n_0_0_157));
   OAI21_X1 i_0_0_163 (.A(n_0_0_159), .B1(n_0_0_178), .B2(\values[6] [4]), 
      .ZN(n_0_0_158));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_178), .A2(n_0_0_213), .ZN(n_0_0_159));
   OAI21_X1 i_0_0_165 (.A(n_0_0_161), .B1(n_0_0_163), .B2(n_0_0_162), .ZN(
      n_0_0_160));
   AOI22_X1 i_0_0_166 (.A1(\values[7] [3]), .A2(n_0_0_171), .B1(n_0_0_169), 
      .B2(\values[7] [2]), .ZN(n_0_0_161));
   OAI22_X1 i_0_0_167 (.A1(\values[7] [2]), .A2(n_0_0_169), .B1(n_0_0_164), 
      .B2(\values[7] [1]), .ZN(n_0_0_162));
   AOI22_X1 i_0_0_168 (.A1(\values[7] [0]), .A2(n_0_0_166), .B1(n_0_0_164), 
      .B2(\values[7] [1]), .ZN(n_0_0_163));
   OAI21_X1 i_0_0_169 (.A(n_0_0_165), .B1(n_0_0_178), .B2(\values[6] [1]), 
      .ZN(n_0_0_164));
   NAND2_X1 i_0_0_170 (.A1(n_0_0_178), .A2(n_0_0_224), .ZN(n_0_0_165));
   INV_X1 i_0_0_171 (.A(n_0_0_167), .ZN(n_0_0_166));
   OAI21_X1 i_0_0_172 (.A(n_0_0_168), .B1(n_0_0_177), .B2(n_0_0_221), .ZN(
      n_0_0_167));
   NAND2_X1 i_0_0_173 (.A1(\values[6] [0]), .A2(n_0_0_177), .ZN(n_0_0_168));
   OAI21_X1 i_0_0_174 (.A(n_0_0_170), .B1(n_0_0_178), .B2(\values[6] [2]), 
      .ZN(n_0_0_169));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_226), .A2(n_0_0_178), .ZN(n_0_0_170));
   OAI21_X1 i_0_0_176 (.A(n_0_0_172), .B1(n_0_0_178), .B2(\values[6] [3]), 
      .ZN(n_0_0_171));
   NAND2_X1 i_0_0_177 (.A1(n_0_0_178), .A2(n_0_0_217), .ZN(n_0_0_172));
   OAI21_X1 i_0_0_178 (.A(n_0_0_174), .B1(n_0_0_178), .B2(\values[6] [8]), 
      .ZN(n_0_0_173));
   NAND2_X1 i_0_0_179 (.A1(n_0_0_200), .A2(n_0_0_178), .ZN(n_0_0_174));
   NAND2_X1 i_0_0_180 (.A1(\values[6] [15]), .A2(n_0_0_236), .ZN(n_0_0_175));
   AND2_X1 i_0_0_181 (.A1(\values[6] [15]), .A2(n_0_0_236), .ZN(n_0_0_176));
   INV_X1 i_0_0_182 (.A(n_0_0_178), .ZN(n_0_0_177));
   OR2_X1 i_0_0_183 (.A1(n_0_0_180), .A2(n_0_0_179), .ZN(n_0_0_178));
   NOR2_X1 i_0_0_184 (.A1(n_0_0_236), .A2(n_0_0_181), .ZN(n_0_0_179));
   AOI21_X1 i_0_0_185 (.A(n_0_0_508), .B1(n_0_0_236), .B2(n_0_0_181), .ZN(
      n_0_0_180));
   OAI21_X1 i_0_0_186 (.A(n_0_0_232), .B1(n_0_0_182), .B2(n_0_0_233), .ZN(
      n_0_0_181));
   OAI21_X1 i_0_0_187 (.A(n_0_0_183), .B1(n_0_0_230), .B2(\values[6] [13]), 
      .ZN(n_0_0_182));
   NAND3_X1 i_0_0_188 (.A1(n_0_0_188), .A2(n_0_0_185), .A3(n_0_0_184), .ZN(
      n_0_0_183));
   NAND2_X1 i_0_0_189 (.A1(n_0_0_230), .A2(\values[6] [13]), .ZN(n_0_0_184));
   OAI221_X1 i_0_0_190 (.A(n_0_0_186), .B1(n_0_0_190), .B2(\values[6] [11]), 
      .C1(\values[6] [12]), .C2(n_0_0_228), .ZN(n_0_0_185));
   OAI21_X1 i_0_0_191 (.A(n_0_0_187), .B1(n_0_0_189), .B2(n_0_0_192), .ZN(
      n_0_0_186));
   NAND2_X1 i_0_0_192 (.A1(n_0_0_190), .A2(\values[6] [11]), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_193 (.A1(n_0_0_228), .A2(\values[6] [12]), .ZN(n_0_0_188));
   NOR2_X1 i_0_0_194 (.A1(n_0_0_193), .A2(\values[6] [10]), .ZN(n_0_0_189));
   AOI21_X1 i_0_0_195 (.A(n_0_0_191), .B1(n_0_0_238), .B2(\values[5] [11]), 
      .ZN(n_0_0_190));
   NOR2_X1 i_0_0_196 (.A1(n_0_0_238), .A2(n_0_0_255), .ZN(n_0_0_191));
   AOI221_X1 i_0_0_197 (.A(n_0_0_195), .B1(n_0_0_193), .B2(\values[6] [10]), 
      .C1(\values[6] [9]), .C2(n_0_0_197), .ZN(n_0_0_192));
   AOI21_X1 i_0_0_198 (.A(n_0_0_194), .B1(n_0_0_238), .B2(\values[5] [10]), 
      .ZN(n_0_0_193));
   NOR2_X1 i_0_0_199 (.A1(n_0_0_238), .A2(n_0_0_258), .ZN(n_0_0_194));
   AOI21_X1 i_0_0_200 (.A(n_0_0_196), .B1(n_0_0_202), .B2(n_0_0_199), .ZN(
      n_0_0_195));
   OAI22_X1 i_0_0_201 (.A1(\values[6] [8]), .A2(n_0_0_200), .B1(n_0_0_197), 
      .B2(\values[6] [9]), .ZN(n_0_0_196));
   AOI21_X1 i_0_0_202 (.A(n_0_0_198), .B1(n_0_0_238), .B2(\values[5] [9]), 
      .ZN(n_0_0_197));
   NOR2_X1 i_0_0_203 (.A1(n_0_0_262), .A2(n_0_0_238), .ZN(n_0_0_198));
   AOI22_X1 i_0_0_204 (.A1(\values[6] [7]), .A2(n_0_0_203), .B1(n_0_0_200), 
      .B2(\values[6] [8]), .ZN(n_0_0_199));
   AOI21_X1 i_0_0_205 (.A(n_0_0_201), .B1(n_0_0_238), .B2(\values[5] [8]), 
      .ZN(n_0_0_200));
   NOR2_X1 i_0_0_206 (.A1(n_0_0_238), .A2(n_0_0_265), .ZN(n_0_0_201));
   OAI221_X1 i_0_0_207 (.A(n_0_0_205), .B1(n_0_0_203), .B2(\values[6] [7]), 
      .C1(\values[6] [6]), .C2(n_0_0_207), .ZN(n_0_0_202));
   AOI21_X1 i_0_0_208 (.A(n_0_0_204), .B1(n_0_0_238), .B2(\values[5] [7]), 
      .ZN(n_0_0_203));
   NOR2_X1 i_0_0_209 (.A1(n_0_0_238), .A2(n_0_0_268), .ZN(n_0_0_204));
   OAI21_X1 i_0_0_210 (.A(n_0_0_206), .B1(n_0_0_212), .B2(n_0_0_209), .ZN(
      n_0_0_205));
   AOI22_X1 i_0_0_211 (.A1(\values[6] [5]), .A2(n_0_0_210), .B1(n_0_0_207), 
      .B2(\values[6] [6]), .ZN(n_0_0_206));
   AOI21_X1 i_0_0_212 (.A(n_0_0_208), .B1(n_0_0_238), .B2(\values[5] [6]), 
      .ZN(n_0_0_207));
   NOR2_X1 i_0_0_213 (.A1(n_0_0_238), .A2(n_0_0_272), .ZN(n_0_0_208));
   OAI22_X1 i_0_0_214 (.A1(\values[6] [4]), .A2(n_0_0_213), .B1(n_0_0_210), 
      .B2(\values[6] [5]), .ZN(n_0_0_209));
   AOI21_X1 i_0_0_215 (.A(n_0_0_211), .B1(n_0_0_238), .B2(\values[5] [5]), 
      .ZN(n_0_0_210));
   NOR2_X1 i_0_0_216 (.A1(n_0_0_238), .A2(n_0_0_275), .ZN(n_0_0_211));
   AOI221_X1 i_0_0_217 (.A(n_0_0_215), .B1(n_0_0_213), .B2(\values[6] [4]), 
      .C1(\values[6] [3]), .C2(n_0_0_217), .ZN(n_0_0_212));
   AOI21_X1 i_0_0_218 (.A(n_0_0_214), .B1(n_0_0_238), .B2(\values[5] [4]), 
      .ZN(n_0_0_213));
   NOR2_X1 i_0_0_219 (.A1(n_0_0_238), .A2(n_0_0_278), .ZN(n_0_0_214));
   AOI21_X1 i_0_0_220 (.A(n_0_0_216), .B1(n_0_0_219), .B2(n_0_0_220), .ZN(
      n_0_0_215));
   OAI22_X1 i_0_0_221 (.A1(\values[6] [2]), .A2(n_0_0_226), .B1(n_0_0_217), 
      .B2(\values[6] [3]), .ZN(n_0_0_216));
   AOI21_X1 i_0_0_222 (.A(n_0_0_218), .B1(n_0_0_238), .B2(\values[5] [3]), 
      .ZN(n_0_0_217));
   NOR2_X1 i_0_0_223 (.A1(n_0_0_238), .A2(n_0_0_282), .ZN(n_0_0_218));
   AOI22_X1 i_0_0_224 (.A1(\values[6] [2]), .A2(n_0_0_226), .B1(n_0_0_224), 
      .B2(\values[6] [1]), .ZN(n_0_0_219));
   OAI211_X1 i_0_0_225 (.A(\values[6] [0]), .B(n_0_0_221), .C1(n_0_0_224), 
      .C2(\values[6] [1]), .ZN(n_0_0_220));
   INV_X1 i_0_0_226 (.A(n_0_0_222), .ZN(n_0_0_221));
   OAI21_X1 i_0_0_227 (.A(n_0_0_223), .B1(n_0_0_238), .B2(n_0_0_290), .ZN(
      n_0_0_222));
   NAND2_X1 i_0_0_228 (.A1(n_0_0_238), .A2(\values[5] [0]), .ZN(n_0_0_223));
   AOI21_X1 i_0_0_229 (.A(n_0_0_225), .B1(n_0_0_238), .B2(\values[5] [1]), 
      .ZN(n_0_0_224));
   NOR2_X1 i_0_0_230 (.A1(n_0_0_238), .A2(n_0_0_288), .ZN(n_0_0_225));
   AOI21_X1 i_0_0_231 (.A(n_0_0_227), .B1(n_0_0_238), .B2(\values[5] [2]), 
      .ZN(n_0_0_226));
   NOR2_X1 i_0_0_232 (.A1(n_0_0_238), .A2(n_0_0_285), .ZN(n_0_0_227));
   AOI21_X1 i_0_0_233 (.A(n_0_0_229), .B1(n_0_0_238), .B2(\values[5] [12]), 
      .ZN(n_0_0_228));
   NOR2_X1 i_0_0_234 (.A1(n_0_0_238), .A2(n_0_0_252), .ZN(n_0_0_229));
   AOI21_X1 i_0_0_235 (.A(n_0_0_231), .B1(n_0_0_238), .B2(\values[5] [13]), 
      .ZN(n_0_0_230));
   NOR2_X1 i_0_0_236 (.A1(n_0_0_248), .A2(n_0_0_238), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_237 (.A1(n_0_0_234), .A2(\values[6] [14]), .ZN(n_0_0_232));
   NOR2_X1 i_0_0_238 (.A1(n_0_0_234), .A2(\values[6] [14]), .ZN(n_0_0_233));
   AOI21_X1 i_0_0_239 (.A(n_0_0_235), .B1(n_0_0_238), .B2(\values[5] [14]), 
      .ZN(n_0_0_234));
   NOR2_X1 i_0_0_240 (.A1(n_0_0_245), .A2(n_0_0_238), .ZN(n_0_0_235));
   NOR2_X1 i_0_0_241 (.A1(n_0_0_509), .A2(n_0_0_243), .ZN(n_0_0_236));
   NOR2_X1 i_0_0_242 (.A1(n_0_0_292), .A2(n_0_0_238), .ZN(n_0_0_237));
   OAI211_X1 i_0_0_243 (.A(n_0_0_240), .B(n_0_0_239), .C1(\values[5] [15]), 
      .C2(n_0_0_243), .ZN(n_0_0_238));
   OAI211_X1 i_0_0_244 (.A(n_0_0_245), .B(\values[5] [14]), .C1(n_0_0_509), 
      .C2(n_0_0_242), .ZN(n_0_0_239));
   OAI21_X1 i_0_0_245 (.A(n_0_0_241), .B1(n_0_0_248), .B2(\values[5] [13]), 
      .ZN(n_0_0_240));
   AOI211_X1 i_0_0_246 (.A(n_0_0_247), .B(n_0_0_244), .C1(n_0_0_243), .C2(
      \values[5] [15]), .ZN(n_0_0_241));
   INV_X1 i_0_0_247 (.A(n_0_0_243), .ZN(n_0_0_242));
   NAND3_X1 i_0_0_248 (.A1(\values[3] [15]), .A2(\values[4] [15]), .A3(n_0_0_359), 
      .ZN(n_0_0_243));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_245), .A2(\values[5] [14]), .ZN(n_0_0_244));
   AOI21_X1 i_0_0_250 (.A(n_0_0_246), .B1(n_0_0_292), .B2(\values[4] [14]), 
      .ZN(n_0_0_245));
   NOR2_X1 i_0_0_251 (.A1(n_0_0_297), .A2(n_0_0_292), .ZN(n_0_0_246));
   AOI221_X1 i_0_0_252 (.A(n_0_0_250), .B1(n_0_0_248), .B2(\values[5] [13]), 
      .C1(\values[5] [12]), .C2(n_0_0_252), .ZN(n_0_0_247));
   AOI21_X1 i_0_0_253 (.A(n_0_0_249), .B1(n_0_0_292), .B2(\values[4] [13]), 
      .ZN(n_0_0_248));
   NOR2_X1 i_0_0_254 (.A1(n_0_0_300), .A2(n_0_0_292), .ZN(n_0_0_249));
   AOI21_X1 i_0_0_255 (.A(n_0_0_251), .B1(n_0_0_257), .B2(n_0_0_254), .ZN(
      n_0_0_250));
   OAI22_X1 i_0_0_256 (.A1(\values[5] [11]), .A2(n_0_0_255), .B1(n_0_0_252), 
      .B2(\values[5] [12]), .ZN(n_0_0_251));
   AOI21_X1 i_0_0_257 (.A(n_0_0_253), .B1(n_0_0_292), .B2(\values[4] [12]), 
      .ZN(n_0_0_252));
   NOR2_X1 i_0_0_258 (.A1(n_0_0_303), .A2(n_0_0_292), .ZN(n_0_0_253));
   AOI22_X1 i_0_0_259 (.A1(\values[5] [10]), .A2(n_0_0_258), .B1(n_0_0_255), 
      .B2(\values[5] [11]), .ZN(n_0_0_254));
   AOI21_X1 i_0_0_260 (.A(n_0_0_256), .B1(n_0_0_292), .B2(\values[4] [11]), 
      .ZN(n_0_0_255));
   NOR2_X1 i_0_0_261 (.A1(n_0_0_307), .A2(n_0_0_292), .ZN(n_0_0_256));
   OAI221_X1 i_0_0_262 (.A(n_0_0_260), .B1(n_0_0_258), .B2(\values[5] [10]), 
      .C1(\values[5] [9]), .C2(n_0_0_262), .ZN(n_0_0_257));
   AOI21_X1 i_0_0_263 (.A(n_0_0_259), .B1(n_0_0_292), .B2(\values[4] [10]), 
      .ZN(n_0_0_258));
   NOR2_X1 i_0_0_264 (.A1(n_0_0_311), .A2(n_0_0_292), .ZN(n_0_0_259));
   OAI21_X1 i_0_0_265 (.A(n_0_0_261), .B1(n_0_0_267), .B2(n_0_0_264), .ZN(
      n_0_0_260));
   AOI22_X1 i_0_0_266 (.A1(\values[5] [8]), .A2(n_0_0_265), .B1(n_0_0_262), 
      .B2(\values[5] [9]), .ZN(n_0_0_261));
   AOI21_X1 i_0_0_267 (.A(n_0_0_263), .B1(n_0_0_292), .B2(\values[4] [9]), 
      .ZN(n_0_0_262));
   NOR2_X1 i_0_0_268 (.A1(n_0_0_314), .A2(n_0_0_292), .ZN(n_0_0_263));
   OAI22_X1 i_0_0_269 (.A1(\values[5] [7]), .A2(n_0_0_268), .B1(n_0_0_265), 
      .B2(\values[5] [8]), .ZN(n_0_0_264));
   AOI21_X1 i_0_0_270 (.A(n_0_0_266), .B1(n_0_0_292), .B2(\values[4] [8]), 
      .ZN(n_0_0_265));
   NOR2_X1 i_0_0_271 (.A1(n_0_0_317), .A2(n_0_0_292), .ZN(n_0_0_266));
   AOI221_X1 i_0_0_272 (.A(n_0_0_270), .B1(n_0_0_268), .B2(\values[5] [7]), 
      .C1(\values[5] [6]), .C2(n_0_0_272), .ZN(n_0_0_267));
   AOI21_X1 i_0_0_273 (.A(n_0_0_269), .B1(n_0_0_292), .B2(\values[4] [7]), 
      .ZN(n_0_0_268));
   NOR2_X1 i_0_0_274 (.A1(n_0_0_321), .A2(n_0_0_292), .ZN(n_0_0_269));
   AOI21_X1 i_0_0_275 (.A(n_0_0_271), .B1(n_0_0_277), .B2(n_0_0_274), .ZN(
      n_0_0_270));
   OAI22_X1 i_0_0_276 (.A1(\values[5] [5]), .A2(n_0_0_275), .B1(n_0_0_272), 
      .B2(\values[5] [6]), .ZN(n_0_0_271));
   AOI21_X1 i_0_0_277 (.A(n_0_0_273), .B1(n_0_0_292), .B2(\values[4] [6]), 
      .ZN(n_0_0_272));
   NOR2_X1 i_0_0_278 (.A1(n_0_0_324), .A2(n_0_0_292), .ZN(n_0_0_273));
   AOI22_X1 i_0_0_279 (.A1(\values[5] [4]), .A2(n_0_0_278), .B1(n_0_0_275), 
      .B2(\values[5] [5]), .ZN(n_0_0_274));
   AOI21_X1 i_0_0_280 (.A(n_0_0_276), .B1(n_0_0_292), .B2(\values[4] [5]), 
      .ZN(n_0_0_275));
   NOR2_X1 i_0_0_281 (.A1(n_0_0_328), .A2(n_0_0_292), .ZN(n_0_0_276));
   OAI221_X1 i_0_0_282 (.A(n_0_0_280), .B1(n_0_0_278), .B2(\values[5] [4]), 
      .C1(\values[5] [3]), .C2(n_0_0_282), .ZN(n_0_0_277));
   AOI21_X1 i_0_0_283 (.A(n_0_0_279), .B1(n_0_0_292), .B2(\values[4] [4]), 
      .ZN(n_0_0_278));
   NOR2_X1 i_0_0_284 (.A1(n_0_0_331), .A2(n_0_0_292), .ZN(n_0_0_279));
   OAI21_X1 i_0_0_285 (.A(n_0_0_281), .B1(n_0_0_287), .B2(n_0_0_284), .ZN(
      n_0_0_280));
   AOI22_X1 i_0_0_286 (.A1(\values[5] [2]), .A2(n_0_0_285), .B1(n_0_0_282), 
      .B2(\values[5] [3]), .ZN(n_0_0_281));
   AOI21_X1 i_0_0_287 (.A(n_0_0_283), .B1(n_0_0_292), .B2(\values[4] [3]), 
      .ZN(n_0_0_282));
   NOR2_X1 i_0_0_288 (.A1(n_0_0_334), .A2(n_0_0_292), .ZN(n_0_0_283));
   OAI22_X1 i_0_0_289 (.A1(\values[5] [1]), .A2(n_0_0_288), .B1(n_0_0_285), 
      .B2(\values[5] [2]), .ZN(n_0_0_284));
   AOI21_X1 i_0_0_290 (.A(n_0_0_286), .B1(n_0_0_292), .B2(\values[4] [2]), 
      .ZN(n_0_0_285));
   NOR2_X1 i_0_0_291 (.A1(n_0_0_338), .A2(n_0_0_292), .ZN(n_0_0_286));
   AOI22_X1 i_0_0_292 (.A1(\values[5] [0]), .A2(n_0_0_290), .B1(n_0_0_288), 
      .B2(\values[5] [1]), .ZN(n_0_0_287));
   OAI21_X1 i_0_0_293 (.A(n_0_0_289), .B1(n_0_0_292), .B2(n_0_0_342), .ZN(
      n_0_0_288));
   NAND2_X1 i_0_0_294 (.A1(n_0_0_510), .A2(n_0_0_292), .ZN(n_0_0_289));
   INV_X1 i_0_0_295 (.A(n_0_0_291), .ZN(n_0_0_290));
   MUX2_X1 i_0_0_296 (.A(n_0_0_341), .B(\values[4] [0]), .S(n_0_0_292), .Z(
      n_0_0_291));
   OAI21_X1 i_0_0_297 (.A(n_0_0_293), .B1(n_0_0_344), .B2(\values[4] [15]), 
      .ZN(n_0_0_292));
   OAI211_X1 i_0_0_298 (.A(n_0_0_295), .B(n_0_0_294), .C1(\values[4] [14]), 
      .C2(n_0_0_297), .ZN(n_0_0_293));
   NAND2_X1 i_0_0_299 (.A1(n_0_0_344), .A2(\values[4] [15]), .ZN(n_0_0_294));
   OAI21_X1 i_0_0_300 (.A(n_0_0_296), .B1(n_0_0_302), .B2(n_0_0_299), .ZN(
      n_0_0_295));
   AOI22_X1 i_0_0_301 (.A1(\values[4] [13]), .A2(n_0_0_300), .B1(n_0_0_297), 
      .B2(\values[4] [14]), .ZN(n_0_0_296));
   OAI21_X1 i_0_0_302 (.A(n_0_0_298), .B1(n_0_0_355), .B2(\values[3] [14]), 
      .ZN(n_0_0_297));
   NAND2_X1 i_0_0_303 (.A1(n_0_0_362), .A2(n_0_0_355), .ZN(n_0_0_298));
   OAI22_X1 i_0_0_304 (.A1(\values[4] [12]), .A2(n_0_0_303), .B1(n_0_0_300), 
      .B2(\values[4] [13]), .ZN(n_0_0_299));
   OAI21_X1 i_0_0_305 (.A(n_0_0_301), .B1(n_0_0_355), .B2(\values[3] [13]), 
      .ZN(n_0_0_300));
   NAND2_X1 i_0_0_306 (.A1(n_0_0_366), .A2(n_0_0_355), .ZN(n_0_0_301));
   AOI222_X1 i_0_0_307 (.A1(n_0_0_309), .A2(n_0_0_305), .B1(n_0_0_303), .B2(
      \values[4] [12]), .C1(\values[4] [11]), .C2(n_0_0_307), .ZN(n_0_0_302));
   OAI21_X1 i_0_0_308 (.A(n_0_0_304), .B1(n_0_0_356), .B2(n_0_0_370), .ZN(
      n_0_0_303));
   NAND2_X1 i_0_0_309 (.A1(n_0_0_356), .A2(n_0_0_511), .ZN(n_0_0_304));
   INV_X1 i_0_0_310 (.A(n_0_0_306), .ZN(n_0_0_305));
   OAI22_X1 i_0_0_311 (.A1(\values[4] [10]), .A2(n_0_0_311), .B1(n_0_0_307), 
      .B2(\values[4] [11]), .ZN(n_0_0_306));
   OAI21_X1 i_0_0_312 (.A(n_0_0_308), .B1(n_0_0_355), .B2(\values[3] [11]), 
      .ZN(n_0_0_307));
   NAND2_X1 i_0_0_313 (.A1(n_0_0_376), .A2(n_0_0_355), .ZN(n_0_0_308));
   OAI21_X1 i_0_0_314 (.A(n_0_0_310), .B1(n_0_0_316), .B2(n_0_0_313), .ZN(
      n_0_0_309));
   AOI22_X1 i_0_0_315 (.A1(\values[4] [9]), .A2(n_0_0_314), .B1(n_0_0_311), 
      .B2(\values[4] [10]), .ZN(n_0_0_310));
   OAI21_X1 i_0_0_316 (.A(n_0_0_312), .B1(n_0_0_355), .B2(\values[3] [10]), 
      .ZN(n_0_0_311));
   NAND2_X1 i_0_0_317 (.A1(n_0_0_379), .A2(n_0_0_355), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_318 (.A1(\values[4] [8]), .A2(n_0_0_317), .B1(n_0_0_314), 
      .B2(\values[4] [9]), .ZN(n_0_0_313));
   AOI21_X1 i_0_0_319 (.A(n_0_0_315), .B1(n_0_0_356), .B2(\values[3] [9]), 
      .ZN(n_0_0_314));
   NOR2_X1 i_0_0_320 (.A1(n_0_0_356), .A2(n_0_0_382), .ZN(n_0_0_315));
   AOI221_X1 i_0_0_321 (.A(n_0_0_319), .B1(n_0_0_317), .B2(\values[4] [8]), 
      .C1(\values[4] [7]), .C2(n_0_0_321), .ZN(n_0_0_316));
   OAI21_X1 i_0_0_322 (.A(n_0_0_318), .B1(n_0_0_355), .B2(\values[3] [8]), 
      .ZN(n_0_0_317));
   NAND2_X1 i_0_0_323 (.A1(n_0_0_387), .A2(n_0_0_355), .ZN(n_0_0_318));
   NOR2_X1 i_0_0_324 (.A1(n_0_0_323), .A2(n_0_0_320), .ZN(n_0_0_319));
   OAI22_X1 i_0_0_325 (.A1(\values[4] [6]), .A2(n_0_0_324), .B1(n_0_0_321), 
      .B2(\values[4] [7]), .ZN(n_0_0_320));
   OAI21_X1 i_0_0_326 (.A(n_0_0_322), .B1(n_0_0_355), .B2(\values[3] [7]), 
      .ZN(n_0_0_321));
   NAND2_X1 i_0_0_327 (.A1(n_0_0_390), .A2(n_0_0_355), .ZN(n_0_0_322));
   AOI221_X1 i_0_0_328 (.A(n_0_0_326), .B1(n_0_0_324), .B2(\values[4] [6]), 
      .C1(\values[4] [5]), .C2(n_0_0_328), .ZN(n_0_0_323));
   OAI21_X1 i_0_0_329 (.A(n_0_0_325), .B1(n_0_0_355), .B2(\values[3] [6]), 
      .ZN(n_0_0_324));
   NAND2_X1 i_0_0_330 (.A1(n_0_0_355), .A2(n_0_0_393), .ZN(n_0_0_325));
   AOI21_X1 i_0_0_331 (.A(n_0_0_327), .B1(n_0_0_333), .B2(n_0_0_330), .ZN(
      n_0_0_326));
   OAI22_X1 i_0_0_332 (.A1(\values[4] [4]), .A2(n_0_0_331), .B1(n_0_0_328), 
      .B2(\values[4] [5]), .ZN(n_0_0_327));
   OAI21_X1 i_0_0_333 (.A(n_0_0_329), .B1(n_0_0_355), .B2(\values[3] [5]), 
      .ZN(n_0_0_328));
   NAND2_X1 i_0_0_334 (.A1(n_0_0_415), .A2(n_0_0_355), .ZN(n_0_0_329));
   AOI22_X1 i_0_0_335 (.A1(\values[4] [3]), .A2(n_0_0_334), .B1(n_0_0_331), 
      .B2(\values[4] [4]), .ZN(n_0_0_330));
   OAI21_X1 i_0_0_336 (.A(n_0_0_332), .B1(n_0_0_355), .B2(\values[3] [4]), 
      .ZN(n_0_0_331));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_412), .A2(n_0_0_355), .ZN(n_0_0_332));
   OAI221_X1 i_0_0_338 (.A(n_0_0_336), .B1(n_0_0_334), .B2(\values[4] [3]), 
      .C1(\values[4] [2]), .C2(n_0_0_338), .ZN(n_0_0_333));
   OAI21_X1 i_0_0_339 (.A(n_0_0_335), .B1(n_0_0_355), .B2(\values[3] [3]), 
      .ZN(n_0_0_334));
   NAND2_X1 i_0_0_340 (.A1(n_0_0_410), .A2(n_0_0_355), .ZN(n_0_0_335));
   OAI21_X1 i_0_0_341 (.A(n_0_0_337), .B1(n_0_0_342), .B2(n_0_0_510), .ZN(
      n_0_0_336));
   AOI22_X1 i_0_0_342 (.A1(\values[4] [0]), .A2(n_0_0_340), .B1(n_0_0_338), 
      .B2(\values[4] [2]), .ZN(n_0_0_337));
   OAI21_X1 i_0_0_343 (.A(n_0_0_339), .B1(n_0_0_355), .B2(\values[3] [2]), 
      .ZN(n_0_0_338));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_402), .A2(n_0_0_355), .ZN(n_0_0_339));
   AOI21_X1 i_0_0_345 (.A(n_0_0_341), .B1(n_0_0_342), .B2(n_0_0_510), .ZN(
      n_0_0_340));
   MUX2_X1 i_0_0_346 (.A(n_0_0_405), .B(\values[3] [0]), .S(n_0_0_356), .Z(
      n_0_0_341));
   OAI21_X1 i_0_0_347 (.A(n_0_0_343), .B1(n_0_0_356), .B2(n_0_0_407), .ZN(
      n_0_0_342));
   NAND2_X1 i_0_0_348 (.A1(\values[3] [1]), .A2(n_0_0_356), .ZN(n_0_0_343));
   NAND2_X1 i_0_0_349 (.A1(\values[3] [15]), .A2(n_0_0_359), .ZN(n_0_0_344));
   INV_X1 i_0_0_350 (.A(n_0_0_346), .ZN(n_0_0_345));
   NOR2_X1 i_0_0_351 (.A1(n_0_0_354), .A2(n_0_0_348), .ZN(n_0_0_346));
   INV_X1 i_0_0_352 (.A(n_0_0_348), .ZN(n_0_0_347));
   NAND2_X1 i_0_0_353 (.A1(n_0_0_478), .A2(n_0_0_349), .ZN(n_0_0_348));
   AND4_X1 i_0_0_354 (.A1(n_0_0_353), .A2(n_0_0_352), .A3(n_0_0_351), .A4(
      n_0_0_350), .ZN(n_0_0_349));
   NOR4_X1 i_0_0_355 (.A1(\values[0] [7]), .A2(\values[0] [6]), .A3(
      \values[0] [5]), .A4(\values[0] [4]), .ZN(n_0_0_350));
   NOR4_X1 i_0_0_356 (.A1(\values[0] [3]), .A2(\values[0] [2]), .A3(
      \values[0] [1]), .A4(\values[0] [0]), .ZN(n_0_0_351));
   NOR4_X1 i_0_0_357 (.A1(n_0_0_526), .A2(\values[0] [14]), .A3(\values[0] [13]), 
      .A4(\values[0] [12]), .ZN(n_0_0_352));
   NOR4_X1 i_0_0_358 (.A1(\values[0] [11]), .A2(\values[0] [10]), .A3(
      \values[0] [9]), .A4(\values[0] [8]), .ZN(n_0_0_353));
   NAND2_X1 i_0_0_359 (.A1(n_0_0_355), .A2(n_0_0_417), .ZN(n_0_0_354));
   INV_X1 i_0_0_360 (.A(n_0_0_356), .ZN(n_0_0_355));
   AOI22_X1 i_0_0_361 (.A1(n_0_0_361), .A2(n_0_0_357), .B1(n_0_0_360), .B2(
      \values[3] [15]), .ZN(n_0_0_356));
   AOI21_X1 i_0_0_362 (.A(n_0_0_358), .B1(n_0_0_362), .B2(\values[3] [14]), 
      .ZN(n_0_0_357));
   NOR2_X1 i_0_0_363 (.A1(n_0_0_360), .A2(\values[3] [15]), .ZN(n_0_0_358));
   INV_X1 i_0_0_364 (.A(n_0_0_360), .ZN(n_0_0_359));
   NAND3_X1 i_0_0_365 (.A1(\values[0] [15]), .A2(\values[1] [15]), .A3(
      \values[2] [15]), .ZN(n_0_0_360));
   OAI221_X1 i_0_0_366 (.A(n_0_0_364), .B1(n_0_0_362), .B2(\values[3] [14]), 
      .C1(\values[3] [13]), .C2(n_0_0_366), .ZN(n_0_0_361));
   OAI21_X1 i_0_0_367 (.A(n_0_0_363), .B1(n_0_0_417), .B2(\values[2] [14]), 
      .ZN(n_0_0_362));
   NAND2_X1 i_0_0_368 (.A1(n_0_0_423), .A2(n_0_0_417), .ZN(n_0_0_363));
   OAI21_X1 i_0_0_369 (.A(n_0_0_365), .B1(n_0_0_368), .B2(n_0_0_373), .ZN(
      n_0_0_364));
   AOI22_X1 i_0_0_370 (.A1(\values[3] [12]), .A2(n_0_0_369), .B1(n_0_0_366), 
      .B2(\values[3] [13]), .ZN(n_0_0_365));
   OAI21_X1 i_0_0_371 (.A(n_0_0_367), .B1(n_0_0_417), .B2(\values[2] [13]), 
      .ZN(n_0_0_366));
   NAND2_X1 i_0_0_372 (.A1(n_0_0_427), .A2(n_0_0_417), .ZN(n_0_0_367));
   NOR2_X1 i_0_0_373 (.A1(n_0_0_369), .A2(\values[3] [12]), .ZN(n_0_0_368));
   OAI21_X1 i_0_0_374 (.A(n_0_0_372), .B1(n_0_0_417), .B2(\values[2] [12]), 
      .ZN(n_0_0_369));
   OAI21_X1 i_0_0_375 (.A(n_0_0_371), .B1(n_0_0_418), .B2(n_0_0_430), .ZN(
      n_0_0_370));
   NAND2_X1 i_0_0_376 (.A1(n_0_0_418), .A2(\values[2] [12]), .ZN(n_0_0_371));
   NAND2_X1 i_0_0_377 (.A1(n_0_0_417), .A2(n_0_0_430), .ZN(n_0_0_372));
   AOI21_X1 i_0_0_378 (.A(n_0_0_374), .B1(n_0_0_376), .B2(\values[3] [11]), 
      .ZN(n_0_0_373));
   AOI21_X1 i_0_0_379 (.A(n_0_0_375), .B1(n_0_0_381), .B2(n_0_0_378), .ZN(
      n_0_0_374));
   OAI22_X1 i_0_0_380 (.A1(\values[3] [10]), .A2(n_0_0_379), .B1(n_0_0_376), 
      .B2(\values[3] [11]), .ZN(n_0_0_375));
   OAI21_X1 i_0_0_381 (.A(n_0_0_377), .B1(n_0_0_417), .B2(\values[2] [11]), 
      .ZN(n_0_0_376));
   NAND2_X1 i_0_0_382 (.A1(n_0_0_433), .A2(n_0_0_417), .ZN(n_0_0_377));
   AOI22_X1 i_0_0_383 (.A1(\values[3] [9]), .A2(n_0_0_382), .B1(n_0_0_379), 
      .B2(\values[3] [10]), .ZN(n_0_0_378));
   OAI21_X1 i_0_0_384 (.A(n_0_0_380), .B1(n_0_0_417), .B2(\values[2] [10]), 
      .ZN(n_0_0_379));
   NAND2_X1 i_0_0_385 (.A1(n_0_0_476), .A2(n_0_0_417), .ZN(n_0_0_380));
   OAI221_X1 i_0_0_386 (.A(n_0_0_385), .B1(n_0_0_382), .B2(\values[3] [9]), 
      .C1(\values[3] [8]), .C2(n_0_0_387), .ZN(n_0_0_381));
   INV_X1 i_0_0_387 (.A(n_0_0_383), .ZN(n_0_0_382));
   OAI21_X1 i_0_0_388 (.A(n_0_0_384), .B1(n_0_0_418), .B2(n_0_0_438), .ZN(
      n_0_0_383));
   NAND2_X1 i_0_0_389 (.A1(n_0_0_418), .A2(\values[2] [9]), .ZN(n_0_0_384));
   OAI21_X1 i_0_0_390 (.A(n_0_0_386), .B1(n_0_0_392), .B2(n_0_0_389), .ZN(
      n_0_0_385));
   AOI22_X1 i_0_0_391 (.A1(\values[3] [7]), .A2(n_0_0_390), .B1(n_0_0_387), 
      .B2(\values[3] [8]), .ZN(n_0_0_386));
   OAI21_X1 i_0_0_392 (.A(n_0_0_388), .B1(n_0_0_417), .B2(\values[2] [8]), 
      .ZN(n_0_0_387));
   NAND2_X1 i_0_0_393 (.A1(n_0_0_473), .A2(n_0_0_417), .ZN(n_0_0_388));
   OAI22_X1 i_0_0_394 (.A1(\values[3] [6]), .A2(n_0_0_393), .B1(n_0_0_390), 
      .B2(\values[3] [7]), .ZN(n_0_0_389));
   OAI21_X1 i_0_0_395 (.A(n_0_0_391), .B1(n_0_0_417), .B2(\values[2] [7]), 
      .ZN(n_0_0_390));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_417), .A2(n_0_0_470), .ZN(n_0_0_391));
   AOI21_X1 i_0_0_397 (.A(n_0_0_395), .B1(n_0_0_393), .B2(\values[3] [6]), 
      .ZN(n_0_0_392));
   OAI21_X1 i_0_0_398 (.A(n_0_0_394), .B1(n_0_0_417), .B2(\values[2] [6]), 
      .ZN(n_0_0_393));
   NAND2_X1 i_0_0_399 (.A1(n_0_0_417), .A2(n_0_0_468), .ZN(n_0_0_394));
   AOI21_X1 i_0_0_400 (.A(n_0_0_414), .B1(n_0_0_397), .B2(n_0_0_396), .ZN(
      n_0_0_395));
   AOI22_X1 i_0_0_401 (.A1(\values[3] [5]), .A2(n_0_0_415), .B1(n_0_0_412), 
      .B2(\values[3] [4]), .ZN(n_0_0_396));
   OAI21_X1 i_0_0_402 (.A(n_0_0_398), .B1(n_0_0_412), .B2(\values[3] [4]), 
      .ZN(n_0_0_397));
   NAND2_X1 i_0_0_403 (.A1(n_0_0_409), .A2(n_0_0_399), .ZN(n_0_0_398));
   OAI221_X1 i_0_0_404 (.A(n_0_0_400), .B1(n_0_0_402), .B2(\values[3] [2]), 
      .C1(\values[3] [3]), .C2(n_0_0_410), .ZN(n_0_0_399));
   OAI21_X1 i_0_0_405 (.A(n_0_0_401), .B1(n_0_0_404), .B2(n_0_0_405), .ZN(
      n_0_0_400));
   AOI22_X1 i_0_0_406 (.A1(\values[3] [1]), .A2(n_0_0_407), .B1(n_0_0_402), 
      .B2(\values[3] [2]), .ZN(n_0_0_401));
   AOI21_X1 i_0_0_407 (.A(n_0_0_403), .B1(n_0_0_418), .B2(\values[2] [2]), 
      .ZN(n_0_0_402));
   NOR2_X1 i_0_0_408 (.A1(n_0_0_418), .A2(n_0_0_459), .ZN(n_0_0_403));
   OAI21_X1 i_0_0_409 (.A(\values[3] [0]), .B1(n_0_0_407), .B2(\values[3] [1]), 
      .ZN(n_0_0_404));
   OAI21_X1 i_0_0_410 (.A(n_0_0_406), .B1(n_0_0_418), .B2(n_0_0_463), .ZN(
      n_0_0_405));
   NAND2_X1 i_0_0_411 (.A1(n_0_0_418), .A2(\values[2] [0]), .ZN(n_0_0_406));
   OAI21_X1 i_0_0_412 (.A(n_0_0_408), .B1(n_0_0_417), .B2(\values[2] [1]), 
      .ZN(n_0_0_407));
   NAND2_X1 i_0_0_413 (.A1(n_0_0_465), .A2(n_0_0_417), .ZN(n_0_0_408));
   NAND2_X1 i_0_0_414 (.A1(n_0_0_410), .A2(\values[3] [3]), .ZN(n_0_0_409));
   OAI21_X1 i_0_0_415 (.A(n_0_0_411), .B1(n_0_0_417), .B2(\values[2] [3]), 
      .ZN(n_0_0_410));
   NAND2_X1 i_0_0_416 (.A1(n_0_0_456), .A2(n_0_0_417), .ZN(n_0_0_411));
   OAI21_X1 i_0_0_417 (.A(n_0_0_413), .B1(n_0_0_417), .B2(\values[2] [4]), 
      .ZN(n_0_0_412));
   NAND2_X1 i_0_0_418 (.A1(n_0_0_451), .A2(n_0_0_417), .ZN(n_0_0_413));
   NOR2_X1 i_0_0_419 (.A1(n_0_0_415), .A2(\values[3] [5]), .ZN(n_0_0_414));
   OAI21_X1 i_0_0_420 (.A(n_0_0_416), .B1(n_0_0_417), .B2(\values[2] [5]), 
      .ZN(n_0_0_415));
   NAND2_X1 i_0_0_421 (.A1(n_0_0_448), .A2(n_0_0_417), .ZN(n_0_0_416));
   INV_X1 i_0_0_422 (.A(n_0_0_418), .ZN(n_0_0_417));
   OAI22_X1 i_0_0_423 (.A1(n_0_0_419), .A2(n_0_0_422), .B1(\values[2] [15]), 
      .B2(n_0_0_421), .ZN(n_0_0_418));
   OAI21_X1 i_0_0_424 (.A(n_0_0_420), .B1(n_0_0_423), .B2(\values[2] [14]), 
      .ZN(n_0_0_419));
   NAND2_X1 i_0_0_425 (.A1(n_0_0_421), .A2(\values[2] [15]), .ZN(n_0_0_420));
   NAND2_X1 i_0_0_426 (.A1(\values[0] [15]), .A2(\values[1] [15]), .ZN(n_0_0_421));
   AOI221_X1 i_0_0_427 (.A(n_0_0_425), .B1(n_0_0_423), .B2(\values[2] [14]), 
      .C1(\values[2] [13]), .C2(n_0_0_427), .ZN(n_0_0_422));
   OAI21_X1 i_0_0_428 (.A(n_0_0_424), .B1(n_0_0_478), .B2(\values[1] [14]), 
      .ZN(n_0_0_423));
   NAND2_X1 i_0_0_429 (.A1(n_0_0_525), .A2(n_0_0_478), .ZN(n_0_0_424));
   AOI21_X1 i_0_0_430 (.A(n_0_0_426), .B1(n_0_0_432), .B2(n_0_0_429), .ZN(
      n_0_0_425));
   OAI22_X1 i_0_0_431 (.A1(\values[2] [12]), .A2(n_0_0_430), .B1(n_0_0_427), 
      .B2(\values[2] [13]), .ZN(n_0_0_426));
   OAI21_X1 i_0_0_432 (.A(n_0_0_428), .B1(n_0_0_478), .B2(\values[1] [13]), 
      .ZN(n_0_0_427));
   NAND2_X1 i_0_0_433 (.A1(n_0_0_524), .A2(n_0_0_478), .ZN(n_0_0_428));
   AOI22_X1 i_0_0_434 (.A1(\values[2] [11]), .A2(n_0_0_433), .B1(n_0_0_430), 
      .B2(\values[2] [12]), .ZN(n_0_0_429));
   OAI21_X1 i_0_0_435 (.A(n_0_0_431), .B1(n_0_0_478), .B2(\values[1] [12]), 
      .ZN(n_0_0_430));
   NAND2_X1 i_0_0_436 (.A1(n_0_0_523), .A2(n_0_0_478), .ZN(n_0_0_431));
   OAI21_X1 i_0_0_437 (.A(n_0_0_435), .B1(n_0_0_433), .B2(\values[2] [11]), 
      .ZN(n_0_0_432));
   OAI21_X1 i_0_0_438 (.A(n_0_0_434), .B1(n_0_0_478), .B2(\values[1] [11]), 
      .ZN(n_0_0_433));
   NAND2_X1 i_0_0_439 (.A1(n_0_0_522), .A2(n_0_0_478), .ZN(n_0_0_434));
   OAI21_X1 i_0_0_440 (.A(n_0_0_475), .B1(n_0_0_437), .B2(n_0_0_436), .ZN(
      n_0_0_435));
   OAI22_X1 i_0_0_441 (.A1(\values[2] [10]), .A2(n_0_0_476), .B1(n_0_0_438), 
      .B2(\values[2] [9]), .ZN(n_0_0_436));
   AOI21_X1 i_0_0_442 (.A(n_0_0_441), .B1(n_0_0_438), .B2(\values[2] [9]), 
      .ZN(n_0_0_437));
   INV_X1 i_0_0_443 (.A(n_0_0_439), .ZN(n_0_0_438));
   OAI21_X1 i_0_0_444 (.A(n_0_0_440), .B1(n_0_0_478), .B2(n_0_0_514), .ZN(
      n_0_0_439));
   NAND2_X1 i_0_0_445 (.A1(n_0_0_478), .A2(\values[0] [9]), .ZN(n_0_0_440));
   AOI21_X1 i_0_0_446 (.A(n_0_0_472), .B1(n_0_0_443), .B2(n_0_0_442), .ZN(
      n_0_0_441));
   AOI22_X1 i_0_0_447 (.A1(\values[2] [8]), .A2(n_0_0_473), .B1(n_0_0_470), 
      .B2(\values[2] [7]), .ZN(n_0_0_442));
   OAI21_X1 i_0_0_448 (.A(n_0_0_444), .B1(n_0_0_470), .B2(\values[2] [7]), 
      .ZN(n_0_0_443));
   NAND2_X1 i_0_0_449 (.A1(n_0_0_467), .A2(n_0_0_445), .ZN(n_0_0_444));
   OAI221_X1 i_0_0_450 (.A(n_0_0_446), .B1(n_0_0_448), .B2(\values[2] [5]), 
      .C1(\values[2] [6]), .C2(n_0_0_468), .ZN(n_0_0_445));
   OAI21_X1 i_0_0_451 (.A(n_0_0_447), .B1(n_0_0_450), .B2(n_0_0_453), .ZN(
      n_0_0_446));
   AOI22_X1 i_0_0_452 (.A1(\values[2] [4]), .A2(n_0_0_451), .B1(n_0_0_448), 
      .B2(\values[2] [5]), .ZN(n_0_0_447));
   OAI21_X1 i_0_0_453 (.A(n_0_0_449), .B1(n_0_0_479), .B2(\values[0] [5]), 
      .ZN(n_0_0_448));
   NAND2_X1 i_0_0_454 (.A1(n_0_0_479), .A2(n_0_0_513), .ZN(n_0_0_449));
   NOR2_X1 i_0_0_455 (.A1(\values[2] [4]), .A2(n_0_0_451), .ZN(n_0_0_450));
   OAI21_X1 i_0_0_456 (.A(n_0_0_452), .B1(n_0_0_478), .B2(\values[1] [4]), 
      .ZN(n_0_0_451));
   NAND2_X1 i_0_0_457 (.A1(n_0_0_517), .A2(n_0_0_478), .ZN(n_0_0_452));
   AOI21_X1 i_0_0_458 (.A(n_0_0_454), .B1(n_0_0_456), .B2(\values[2] [3]), 
      .ZN(n_0_0_453));
   AOI21_X1 i_0_0_459 (.A(n_0_0_455), .B1(n_0_0_462), .B2(n_0_0_458), .ZN(
      n_0_0_454));
   OAI22_X1 i_0_0_460 (.A1(\values[2] [2]), .A2(n_0_0_459), .B1(n_0_0_456), 
      .B2(\values[2] [3]), .ZN(n_0_0_455));
   OAI21_X1 i_0_0_461 (.A(n_0_0_457), .B1(n_0_0_478), .B2(\values[1] [3]), 
      .ZN(n_0_0_456));
   NAND2_X1 i_0_0_462 (.A1(n_0_0_516), .A2(n_0_0_478), .ZN(n_0_0_457));
   AOI22_X1 i_0_0_463 (.A1(\values[2] [1]), .A2(n_0_0_465), .B1(n_0_0_459), 
      .B2(\values[2] [2]), .ZN(n_0_0_458));
   INV_X1 i_0_0_464 (.A(n_0_0_460), .ZN(n_0_0_459));
   OAI21_X1 i_0_0_465 (.A(n_0_0_461), .B1(n_0_0_478), .B2(n_0_0_512), .ZN(
      n_0_0_460));
   NAND2_X1 i_0_0_466 (.A1(n_0_0_478), .A2(\values[0] [2]), .ZN(n_0_0_461));
   OAI211_X1 i_0_0_467 (.A(n_0_0_463), .B(\values[2] [0]), .C1(\values[2] [1]), 
      .C2(n_0_0_465), .ZN(n_0_0_462));
   INV_X1 i_0_0_468 (.A(n_0_0_464), .ZN(n_0_0_463));
   MUX2_X1 i_0_0_469 (.A(\values[0] [0]), .B(\values[1] [0]), .S(n_0_0_479), 
      .Z(n_0_0_464));
   OAI21_X1 i_0_0_470 (.A(n_0_0_466), .B1(n_0_0_478), .B2(\values[1] [1]), 
      .ZN(n_0_0_465));
   NAND2_X1 i_0_0_471 (.A1(n_0_0_515), .A2(n_0_0_478), .ZN(n_0_0_466));
   NAND2_X1 i_0_0_472 (.A1(n_0_0_468), .A2(\values[2] [6]), .ZN(n_0_0_467));
   OAI21_X1 i_0_0_473 (.A(n_0_0_469), .B1(n_0_0_478), .B2(\values[1] [6]), 
      .ZN(n_0_0_468));
   NAND2_X1 i_0_0_474 (.A1(n_0_0_518), .A2(n_0_0_478), .ZN(n_0_0_469));
   OAI21_X1 i_0_0_475 (.A(n_0_0_471), .B1(n_0_0_478), .B2(\values[1] [7]), 
      .ZN(n_0_0_470));
   NAND2_X1 i_0_0_476 (.A1(n_0_0_519), .A2(n_0_0_478), .ZN(n_0_0_471));
   NOR2_X1 i_0_0_477 (.A1(\values[2] [8]), .A2(n_0_0_473), .ZN(n_0_0_472));
   OAI21_X1 i_0_0_478 (.A(n_0_0_474), .B1(n_0_0_478), .B2(\values[1] [8]), 
      .ZN(n_0_0_473));
   NAND2_X1 i_0_0_479 (.A1(n_0_0_520), .A2(n_0_0_478), .ZN(n_0_0_474));
   NAND2_X1 i_0_0_480 (.A1(\values[2] [10]), .A2(n_0_0_476), .ZN(n_0_0_475));
   OAI21_X1 i_0_0_481 (.A(n_0_0_477), .B1(n_0_0_478), .B2(\values[1] [10]), 
      .ZN(n_0_0_476));
   NAND2_X1 i_0_0_482 (.A1(n_0_0_521), .A2(n_0_0_478), .ZN(n_0_0_477));
   INV_X1 i_0_0_483 (.A(n_0_0_479), .ZN(n_0_0_478));
   AOI21_X1 i_0_0_484 (.A(n_0_0_480), .B1(\values[1] [15]), .B2(n_0_0_526), 
      .ZN(n_0_0_479));
   AOI211_X1 i_0_0_485 (.A(n_0_0_482), .B(n_0_0_481), .C1(n_0_0_525), .C2(
      \values[1] [14]), .ZN(n_0_0_480));
   NOR2_X1 i_0_0_486 (.A1(n_0_0_526), .A2(\values[1] [15]), .ZN(n_0_0_481));
   AOI21_X1 i_0_0_487 (.A(n_0_0_483), .B1(n_0_0_485), .B2(n_0_0_484), .ZN(
      n_0_0_482));
   OAI22_X1 i_0_0_488 (.A1(n_0_0_525), .A2(\values[1] [14]), .B1(n_0_0_524), 
      .B2(\values[1] [13]), .ZN(n_0_0_483));
   AOI22_X1 i_0_0_489 (.A1(n_0_0_524), .A2(\values[1] [13]), .B1(n_0_0_523), 
      .B2(\values[1] [12]), .ZN(n_0_0_484));
   OAI21_X1 i_0_0_490 (.A(n_0_0_486), .B1(\values[1] [11]), .B2(n_0_0_522), 
      .ZN(n_0_0_485));
   AOI21_X1 i_0_0_491 (.A(n_0_0_487), .B1(n_0_0_489), .B2(n_0_0_488), .ZN(
      n_0_0_486));
   NOR2_X1 i_0_0_492 (.A1(n_0_0_523), .A2(\values[1] [12]), .ZN(n_0_0_487));
   AOI22_X1 i_0_0_493 (.A1(n_0_0_522), .A2(\values[1] [11]), .B1(n_0_0_521), 
      .B2(\values[1] [10]), .ZN(n_0_0_488));
   OAI211_X1 i_0_0_494 (.A(n_0_0_491), .B(n_0_0_490), .C1(n_0_0_521), .C2(
      \values[1] [10]), .ZN(n_0_0_489));
   NAND2_X1 i_0_0_495 (.A1(n_0_0_514), .A2(\values[0] [9]), .ZN(n_0_0_490));
   OAI211_X1 i_0_0_496 (.A(n_0_0_493), .B(n_0_0_492), .C1(\values[0] [9]), 
      .C2(n_0_0_514), .ZN(n_0_0_491));
   NAND2_X1 i_0_0_497 (.A1(n_0_0_520), .A2(\values[1] [8]), .ZN(n_0_0_492));
   OAI221_X1 i_0_0_498 (.A(n_0_0_494), .B1(\values[1] [7]), .B2(n_0_0_519), 
      .C1(n_0_0_520), .C2(\values[1] [8]), .ZN(n_0_0_493));
   NAND2_X1 i_0_0_499 (.A1(n_0_0_496), .A2(n_0_0_495), .ZN(n_0_0_494));
   AOI22_X1 i_0_0_500 (.A1(n_0_0_519), .A2(\values[1] [7]), .B1(n_0_0_518), 
      .B2(\values[1] [6]), .ZN(n_0_0_495));
   OAI22_X1 i_0_0_501 (.A1(n_0_0_505), .A2(n_0_0_497), .B1(n_0_0_518), .B2(
      \values[1] [6]), .ZN(n_0_0_496));
   AOI221_X1 i_0_0_502 (.A(n_0_0_498), .B1(n_0_0_513), .B2(\values[0] [5]), 
      .C1(n_0_0_500), .C2(n_0_0_499), .ZN(n_0_0_497));
   NOR2_X1 i_0_0_503 (.A1(n_0_0_517), .A2(\values[1] [4]), .ZN(n_0_0_498));
   AOI22_X1 i_0_0_504 (.A1(n_0_0_517), .A2(\values[1] [4]), .B1(n_0_0_516), 
      .B2(\values[1] [3]), .ZN(n_0_0_499));
   OAI211_X1 i_0_0_505 (.A(n_0_0_502), .B(n_0_0_501), .C1(n_0_0_516), .C2(
      \values[1] [3]), .ZN(n_0_0_500));
   NAND2_X1 i_0_0_506 (.A1(n_0_0_512), .A2(\values[0] [2]), .ZN(n_0_0_501));
   OAI221_X1 i_0_0_507 (.A(n_0_0_503), .B1(\values[0] [2]), .B2(n_0_0_512), 
      .C1(n_0_0_504), .C2(\values[0] [0]), .ZN(n_0_0_502));
   NAND2_X1 i_0_0_508 (.A1(n_0_0_515), .A2(\values[1] [1]), .ZN(n_0_0_503));
   OAI21_X1 i_0_0_509 (.A(\values[1] [0]), .B1(n_0_0_515), .B2(\values[1] [1]), 
      .ZN(n_0_0_504));
   NOR2_X1 i_0_0_510 (.A1(n_0_0_513), .A2(\values[0] [5]), .ZN(n_0_0_505));
   INV_X1 i_0_0_511 (.A(\values[8] [0]), .ZN(n_0_0_506));
   INV_X1 i_0_0_512 (.A(\values[8] [1]), .ZN(n_0_0_507));
   INV_X1 i_0_0_513 (.A(\values[6] [15]), .ZN(n_0_0_508));
   INV_X1 i_0_0_514 (.A(\values[5] [15]), .ZN(n_0_0_509));
   INV_X1 i_0_0_515 (.A(\values[4] [1]), .ZN(n_0_0_510));
   INV_X1 i_0_0_516 (.A(\values[3] [12]), .ZN(n_0_0_511));
   INV_X1 i_0_0_517 (.A(\values[1] [2]), .ZN(n_0_0_512));
   INV_X1 i_0_0_518 (.A(\values[1] [5]), .ZN(n_0_0_513));
   INV_X1 i_0_0_519 (.A(\values[1] [9]), .ZN(n_0_0_514));
   INV_X1 i_0_0_520 (.A(\values[0] [1]), .ZN(n_0_0_515));
   INV_X1 i_0_0_521 (.A(\values[0] [3]), .ZN(n_0_0_516));
   INV_X1 i_0_0_522 (.A(\values[0] [4]), .ZN(n_0_0_517));
   INV_X1 i_0_0_523 (.A(\values[0] [6]), .ZN(n_0_0_518));
   INV_X1 i_0_0_524 (.A(\values[0] [7]), .ZN(n_0_0_519));
   INV_X1 i_0_0_525 (.A(\values[0] [8]), .ZN(n_0_0_520));
   INV_X1 i_0_0_526 (.A(\values[0] [10]), .ZN(n_0_0_521));
   INV_X1 i_0_0_527 (.A(\values[0] [11]), .ZN(n_0_0_522));
   INV_X1 i_0_0_528 (.A(\values[0] [12]), .ZN(n_0_0_523));
   INV_X1 i_0_0_529 (.A(\values[0] [13]), .ZN(n_0_0_524));
   INV_X1 i_0_0_530 (.A(\values[0] [14]), .ZN(n_0_0_525));
   INV_X1 i_0_0_531 (.A(\values[0] [15]), .ZN(n_0_0_526));
endmodule
