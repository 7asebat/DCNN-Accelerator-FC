/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 19:12:47 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2112004273 */

module datapath(\sums[0] , \sums[2] , \r_values[0] , \r_weights[0] , 
      \r_values[1] , \r_weights[1] );
   input [26:0]\sums[0] ;
   output [26:0]\sums[2] ;
   input [15:0]\r_values[0] ;
   input [15:0]\r_weights[0] ;
   input [15:0]\r_values[1] ;
   input [15:0]\r_weights[1] ;

   HA_X1 i_513 (.A(n_495), .B(n_508), .CO(n_514), .S(n_513));
   FA_X1 i_536 (.A(n_502), .B(n_530), .CI(n_524), .CO(n_538), .S(n_537));
   HA_X1 i_537 (.A(n_517), .B(n_514), .CO(n_540), .S(n_539));
   FA_X1 i_567 (.A(n_531), .B(n_557), .CI(n_550), .CO(n_571), .S(n_570));
   FA_X1 i_568 (.A(n_543), .B(n_564), .CI(n_540), .CO(n_573), .S(n_572));
   HA_X1 i_569 (.A(n_538), .B(n_570), .CO(n_575), .S(n_574));
   FA_X1 i_598 (.A(n_558), .B(n_551), .CI(n_544), .CO(n_605), .S(n_604));
   FA_X1 i_599 (.A(n_565), .B(n_599), .CI(n_592), .CO(n_607), .S(n_606));
   FA_X1 i_600 (.A(n_585), .B(n_578), .CI(n_604), .CO(n_609), .S(n_608));
   FA_X1 i_601 (.A(n_571), .B(n_573), .CI(n_608), .CO(n_611), .S(n_610));
   HA_X1 i_602 (.A(n_606), .B(n_575), .CO(n_613), .S(n_612));
   FA_X1 i_639 (.A(n_593), .B(n_586), .CI(n_579), .CO(n_651), .S(n_650));
   FA_X1 i_640 (.A(n_605), .B(n_643), .CI(n_637), .CO(n_653), .S(n_652));
   FA_X1 i_641 (.A(n_630), .B(n_623), .CI(n_616), .CO(n_655), .S(n_654));
   FA_X1 i_642 (.A(n_650), .B(n_607), .CI(n_609), .CO(n_657), .S(n_656));
   FA_X1 i_643 (.A(n_654), .B(n_652), .CI(n_656), .CO(n_659), .S(n_658));
   HA_X1 i_644 (.A(n_613), .B(n_611), .CO(n_661), .S(n_660));
   FA_X1 i_688 (.A(n_624), .B(n_617), .CI(n_651), .CO(n_706), .S(n_705));
   FA_X1 i_689 (.A(n_644), .B(n_692), .CI(n_685), .CO(n_708), .S(n_707));
   FA_X1 i_690 (.A(n_678), .B(n_671), .CI(n_664), .CO(n_710), .S(n_709));
   FA_X1 i_691 (.A(n_705), .B(n_699), .CI(n_655), .CO(n_712), .S(n_711));
   FA_X1 i_692 (.A(n_653), .B(n_709), .CI(n_707), .CO(n_714), .S(n_713));
   FA_X1 i_693 (.A(n_657), .B(n_711), .CI(n_661), .CO(n_716), .S(n_715));
   HA_X1 i_694 (.A(n_659), .B(n_713), .CO(n_718), .S(n_717));
   FA_X1 i_737 (.A(n_693), .B(n_686), .CI(n_679), .CO(n_762), .S(n_761));
   FA_X1 i_738 (.A(n_672), .B(n_665), .CI(n_700), .CO(n_764), .S(n_763));
   FA_X1 i_739 (.A(n_756), .B(n_749), .CI(n_742), .CO(n_766), .S(n_765));
   FA_X1 i_740 (.A(n_735), .B(n_728), .CI(n_721), .CO(n_768), .S(n_767));
   FA_X1 i_741 (.A(n_706), .B(n_763), .CI(n_761), .CO(n_770), .S(n_769));
   FA_X1 i_742 (.A(n_710), .B(n_708), .CI(n_712), .CO(n_772), .S(n_771));
   FA_X1 i_743 (.A(n_767), .B(n_765), .CI(n_771), .CO(n_774), .S(n_773));
   FA_X1 i_744 (.A(n_769), .B(n_714), .CI(n_716), .CO(n_776), .S(n_775));
   HA_X1 i_745 (.A(n_773), .B(n_718), .CO(n_778), .S(n_777));
   FA_X1 i_796 (.A(n_750), .B(n_743), .CI(n_736), .CO(n_830), .S(n_829));
   FA_X1 i_797 (.A(n_729), .B(n_722), .CI(n_762), .CO(n_832), .S(n_831));
   FA_X1 i_798 (.A(n_822), .B(n_816), .CI(n_809), .CO(n_834), .S(n_833));
   FA_X1 i_799 (.A(n_802), .B(n_795), .CI(n_788), .CO(n_836), .S(n_835));
   FA_X1 i_800 (.A(n_781), .B(n_764), .CI(n_831), .CO(n_838), .S(n_837));
   FA_X1 i_801 (.A(n_829), .B(n_768), .CI(n_766), .CO(n_840), .S(n_839));
   FA_X1 i_802 (.A(n_770), .B(n_835), .CI(n_833), .CO(n_842), .S(n_841));
   FA_X1 i_803 (.A(n_837), .B(n_772), .CI(n_839), .CO(n_844), .S(n_843));
   FA_X1 i_804 (.A(n_774), .B(n_841), .CI(n_843), .CO(n_846), .S(n_845));
   HA_X1 i_805 (.A(n_776), .B(n_778), .CO(n_848), .S(n_847));
   FA_X1 i_863 (.A(n_803), .B(n_796), .CI(n_789), .CO(n_907), .S(n_906));
   FA_X1 i_864 (.A(n_782), .B(n_830), .CI(n_823), .CO(n_909), .S(n_908));
   FA_X1 i_865 (.A(n_893), .B(n_886), .CI(n_879), .CO(n_911), .S(n_910));
   FA_X1 i_866 (.A(n_872), .B(n_865), .CI(n_858), .CO(n_913), .S(n_912));
   FA_X1 i_867 (.A(n_851), .B(n_832), .CI(n_906), .CO(n_915), .S(n_914));
   FA_X1 i_868 (.A(n_900), .B(n_836), .CI(n_834), .CO(n_917), .S(n_916));
   FA_X1 i_869 (.A(n_908), .B(n_840), .CI(n_838), .CO(n_919), .S(n_918));
   FA_X1 i_870 (.A(n_912), .B(n_910), .CI(n_914), .CO(n_921), .S(n_920));
   FA_X1 i_871 (.A(n_916), .B(n_842), .CI(n_918), .CO(n_923), .S(n_922));
   FA_X1 i_872 (.A(n_844), .B(n_920), .CI(n_922), .CO(n_925), .S(n_924));
   HA_X1 i_873 (.A(n_846), .B(n_848), .CO(n_927), .S(n_926));
   FA_X1 i_930 (.A(\sums[0] [11]), .B(n_894), .CI(n_887), .CO(n_985), .S(n_984));
   FA_X1 i_931 (.A(n_880), .B(n_873), .CI(n_866), .CO(n_987), .S(n_986));
   FA_X1 i_932 (.A(n_859), .B(n_852), .CI(n_907), .CO(n_989), .S(n_988));
   FA_X1 i_933 (.A(n_901), .B(n_979), .CI(n_972), .CO(n_991), .S(n_990));
   FA_X1 i_934 (.A(n_965), .B(n_958), .CI(n_951), .CO(n_993), .S(n_992));
   FA_X1 i_935 (.A(n_944), .B(n_937), .CI(n_930), .CO(n_995), .S(n_994));
   FA_X1 i_936 (.A(n_909), .B(n_988), .CI(n_986), .CO(n_997), .S(n_996));
   FA_X1 i_937 (.A(n_984), .B(n_913), .CI(n_911), .CO(n_999), .S(n_998));
   FA_X1 i_938 (.A(n_917), .B(n_915), .CI(n_994), .CO(n_1001), .S(n_1000));
   FA_X1 i_939 (.A(n_992), .B(n_990), .CI(n_919), .CO(n_1003), .S(n_1002));
   FA_X1 i_940 (.A(n_998), .B(n_996), .CI(n_921), .CO(n_1005), .S(n_1004));
   FA_X1 i_941 (.A(n_1000), .B(n_1002), .CI(n_923), .CO(n_1007), .S(n_1006));
   FA_X1 i_942 (.A(n_1004), .B(n_927), .CI(n_925), .CO(n_1009), .S(n_1008));
   FA_X1 i_1007 (.A(n_980), .B(n_973), .CI(n_966), .CO(n_1075), .S(n_1074));
   FA_X1 i_1008 (.A(n_959), .B(n_952), .CI(n_945), .CO(n_1077), .S(n_1076));
   FA_X1 i_1009 (.A(n_938), .B(n_931), .CI(n_987), .CO(n_1079), .S(n_1078));
   FA_X1 i_1010 (.A(n_985), .B(n_1067), .CI(n_1061), .CO(n_1081), .S(n_1080));
   FA_X1 i_1011 (.A(n_1054), .B(n_1047), .CI(n_1040), .CO(n_1083), .S(n_1082));
   FA_X1 i_1012 (.A(n_1033), .B(n_1026), .CI(n_1019), .CO(n_1085), .S(n_1084));
   FA_X1 i_1013 (.A(n_1012), .B(n_989), .CI(n_1078), .CO(n_1087), .S(n_1086));
   FA_X1 i_1014 (.A(n_1076), .B(n_1074), .CI(n_995), .CO(n_1089), .S(n_1088));
   FA_X1 i_1015 (.A(n_993), .B(n_991), .CI(n_999), .CO(n_1091), .S(n_1090));
   FA_X1 i_1016 (.A(n_997), .B(n_1084), .CI(n_1082), .CO(n_1093), .S(n_1092));
   FA_X1 i_1017 (.A(n_1080), .B(n_1086), .CI(n_1090), .CO(n_1095), .S(n_1094));
   FA_X1 i_1018 (.A(n_1088), .B(n_1001), .CI(n_1003), .CO(n_1097), .S(n_1096));
   FA_X1 i_1019 (.A(n_1005), .B(n_1092), .CI(n_1094), .CO(n_1099), .S(n_1098));
   FA_X1 i_1020 (.A(n_1096), .B(n_1007), .CI(n_1098), .CO(n_1101), .S(n_1100));
   FA_X1 i_1092 (.A(n_1062), .B(n_1055), .CI(n_1048), .CO(n_1174), .S(n_1173));
   FA_X1 i_1093 (.A(n_1041), .B(n_1034), .CI(n_1027), .CO(n_1176), .S(n_1175));
   FA_X1 i_1094 (.A(n_1020), .B(n_1013), .CI(n_1077), .CO(n_1178), .S(n_1177));
   FA_X1 i_1095 (.A(n_1075), .B(n_1167), .CI(n_1160), .CO(n_1180), .S(n_1179));
   FA_X1 i_1096 (.A(n_1153), .B(n_1146), .CI(n_1139), .CO(n_1182), .S(n_1181));
   FA_X1 i_1097 (.A(n_1132), .B(n_1125), .CI(n_1118), .CO(n_1184), .S(n_1183));
   FA_X1 i_1098 (.A(n_1111), .B(n_1104), .CI(n_1079), .CO(n_1186), .S(n_1185));
   FA_X1 i_1099 (.A(n_1177), .B(n_1175), .CI(n_1173), .CO(n_1188), .S(n_1187));
   FA_X1 i_1100 (.A(n_1085), .B(n_1083), .CI(n_1081), .CO(n_1190), .S(n_1189));
   FA_X1 i_1101 (.A(n_1089), .B(n_1087), .CI(n_1185), .CO(n_1192), .S(n_1191));
   FA_X1 i_1102 (.A(n_1183), .B(n_1181), .CI(n_1179), .CO(n_1194), .S(n_1193));
   FA_X1 i_1103 (.A(n_1091), .B(n_1189), .CI(n_1187), .CO(n_1196), .S(n_1195));
   FA_X1 i_1104 (.A(n_1093), .B(n_1191), .CI(n_1095), .CO(n_1198), .S(n_1197));
   FA_X1 i_1105 (.A(n_1097), .B(n_1193), .CI(n_1195), .CO(n_1200), .S(n_1199));
   FA_X1 i_1106 (.A(n_1099), .B(n_1197), .CI(n_1199), .CO(n_1202), .S(n_1201));
   FA_X1 i_1177 (.A(\sums[0] [14]), .B(n_1161), .CI(n_1154), .CO(n_1274), 
      .S(n_1273));
   FA_X1 i_1178 (.A(n_1147), .B(n_1140), .CI(n_1133), .CO(n_1276), .S(n_1275));
   FA_X1 i_1179 (.A(n_1126), .B(n_1119), .CI(n_1112), .CO(n_1278), .S(n_1277));
   FA_X1 i_1180 (.A(n_1105), .B(n_1176), .CI(n_1174), .CO(n_1280), .S(n_1279));
   FA_X1 i_1181 (.A(n_1168), .B(n_1268), .CI(n_1261), .CO(n_1282), .S(n_1281));
   FA_X1 i_1182 (.A(n_1254), .B(n_1247), .CI(n_1240), .CO(n_1284), .S(n_1283));
   FA_X1 i_1183 (.A(n_1233), .B(n_1226), .CI(n_1219), .CO(n_1286), .S(n_1285));
   FA_X1 i_1184 (.A(n_1212), .B(n_1205), .CI(n_1178), .CO(n_1288), .S(n_1287));
   FA_X1 i_1185 (.A(n_1277), .B(n_1275), .CI(n_1273), .CO(n_1290), .S(n_1289));
   FA_X1 i_1186 (.A(n_1184), .B(n_1182), .CI(n_1180), .CO(n_1292), .S(n_1291));
   FA_X1 i_1187 (.A(n_1186), .B(n_1279), .CI(n_1190), .CO(n_1294), .S(n_1293));
   FA_X1 i_1188 (.A(n_1188), .B(n_1287), .CI(n_1285), .CO(n_1296), .S(n_1295));
   FA_X1 i_1189 (.A(n_1283), .B(n_1281), .CI(n_1291), .CO(n_1298), .S(n_1297));
   FA_X1 i_1190 (.A(n_1289), .B(n_1194), .CI(n_1192), .CO(n_1300), .S(n_1299));
   FA_X1 i_1191 (.A(n_1293), .B(n_1196), .CI(n_1297), .CO(n_1302), .S(n_1301));
   FA_X1 i_1192 (.A(n_1295), .B(n_1198), .CI(n_1299), .CO(n_1304), .S(n_1303));
   FA_X1 i_1193 (.A(n_1301), .B(n_1200), .CI(n_1303), .CO(n_1306), .S(n_1305));
   FA_X1 i_1272 (.A(n_1269), .B(n_1262), .CI(n_1255), .CO(n_1386), .S(n_1385));
   FA_X1 i_1273 (.A(n_1248), .B(n_1241), .CI(n_1234), .CO(n_1388), .S(n_1387));
   FA_X1 i_1274 (.A(n_1227), .B(n_1220), .CI(n_1213), .CO(n_1390), .S(n_1389));
   FA_X1 i_1275 (.A(n_1206), .B(n_1278), .CI(n_1276), .CO(n_1392), .S(n_1391));
   FA_X1 i_1276 (.A(n_1274), .B(n_1378), .CI(n_1372), .CO(n_1394), .S(n_1393));
   FA_X1 i_1277 (.A(n_1365), .B(n_1358), .CI(n_1351), .CO(n_1396), .S(n_1395));
   FA_X1 i_1278 (.A(n_1344), .B(n_1337), .CI(n_1330), .CO(n_1398), .S(n_1397));
   FA_X1 i_1279 (.A(n_1323), .B(n_1316), .CI(n_1309), .CO(n_1400), .S(n_1399));
   FA_X1 i_1280 (.A(n_1280), .B(n_1389), .CI(n_1387), .CO(n_1402), .S(n_1401));
   FA_X1 i_1281 (.A(n_1385), .B(n_1286), .CI(n_1284), .CO(n_1404), .S(n_1403));
   FA_X1 i_1282 (.A(n_1282), .B(n_1288), .CI(n_1391), .CO(n_1406), .S(n_1405));
   FA_X1 i_1283 (.A(n_1292), .B(n_1290), .CI(n_1399), .CO(n_1408), .S(n_1407));
   FA_X1 i_1284 (.A(n_1397), .B(n_1395), .CI(n_1393), .CO(n_1410), .S(n_1409));
   FA_X1 i_1285 (.A(n_1294), .B(n_1403), .CI(n_1401), .CO(n_1412), .S(n_1411));
   FA_X1 i_1286 (.A(n_1296), .B(n_1405), .CI(n_1407), .CO(n_1414), .S(n_1413));
   FA_X1 i_1287 (.A(n_1300), .B(n_1298), .CI(n_1409), .CO(n_1416), .S(n_1415));
   FA_X1 i_1288 (.A(n_1411), .B(n_1302), .CI(n_1413), .CO(n_1418), .S(n_1417));
   FA_X1 i_1289 (.A(n_1415), .B(n_1304), .CI(n_1417), .CO(n_1420), .S(n_1419));
   FA_X1 i_1360 (.A(\sums[0] [16]), .B(n_1379), .CI(n_1373), .CO(n_1492), 
      .S(n_1491));
   FA_X1 i_1361 (.A(n_1366), .B(n_1359), .CI(n_1352), .CO(n_1494), .S(n_1493));
   FA_X1 i_1362 (.A(n_1345), .B(n_1338), .CI(n_1331), .CO(n_1496), .S(n_1495));
   FA_X1 i_1363 (.A(n_1324), .B(n_1317), .CI(n_1310), .CO(n_1498), .S(n_1497));
   FA_X1 i_1364 (.A(n_1390), .B(n_1388), .CI(n_1386), .CO(n_1500), .S(n_1499));
   FA_X1 i_1365 (.A(n_1486), .B(n_1479), .CI(n_1472), .CO(n_1502), .S(n_1501));
   FA_X1 i_1366 (.A(n_1465), .B(n_1458), .CI(n_1451), .CO(n_1504), .S(n_1503));
   FA_X1 i_1367 (.A(n_1444), .B(n_1437), .CI(n_1430), .CO(n_1506), .S(n_1505));
   FA_X1 i_1368 (.A(n_1423), .B(n_1392), .CI(n_1497), .CO(n_1508), .S(n_1507));
   FA_X1 i_1369 (.A(n_1495), .B(n_1493), .CI(n_1491), .CO(n_1510), .S(n_1509));
   FA_X1 i_1370 (.A(n_1400), .B(n_1398), .CI(n_1396), .CO(n_1512), .S(n_1511));
   FA_X1 i_1371 (.A(n_1394), .B(n_1499), .CI(n_1404), .CO(n_1514), .S(n_1513));
   FA_X1 i_1372 (.A(n_1402), .B(n_1505), .CI(n_1503), .CO(n_1516), .S(n_1515));
   FA_X1 i_1373 (.A(n_1501), .B(n_1507), .CI(n_1406), .CO(n_1518), .S(n_1517));
   FA_X1 i_1374 (.A(n_1511), .B(n_1509), .CI(n_1410), .CO(n_1520), .S(n_1519));
   FA_X1 i_1375 (.A(n_1408), .B(n_1513), .CI(n_1412), .CO(n_1522), .S(n_1521));
   FA_X1 i_1376 (.A(n_1515), .B(n_1517), .CI(n_1414), .CO(n_1524), .S(n_1523));
   FA_X1 i_1377 (.A(n_1519), .B(n_1416), .CI(n_1521), .CO(n_1526), .S(n_1525));
   FA_X1 i_1378 (.A(n_1418), .B(n_1523), .CI(n_1525), .CO(n_1528), .S(n_1527));
   FA_X1 i_1450 (.A(n_1480), .B(n_1473), .CI(n_1466), .CO(n_1601), .S(n_1600));
   FA_X1 i_1451 (.A(n_1459), .B(n_1452), .CI(n_1445), .CO(n_1603), .S(n_1602));
   FA_X1 i_1452 (.A(n_1438), .B(n_1431), .CI(n_1424), .CO(n_1605), .S(n_1604));
   FA_X1 i_1453 (.A(n_1498), .B(n_1496), .CI(n_1494), .CO(n_1607), .S(n_1606));
   FA_X1 i_1454 (.A(n_1492), .B(n_1594), .CI(n_1587), .CO(n_1609), .S(n_1608));
   FA_X1 i_1455 (.A(n_1580), .B(n_1573), .CI(n_1566), .CO(n_1611), .S(n_1610));
   FA_X1 i_1456 (.A(n_1559), .B(n_1552), .CI(n_1545), .CO(n_1613), .S(n_1612));
   FA_X1 i_1457 (.A(n_1538), .B(n_1531), .CI(n_1500), .CO(n_1615), .S(n_1614));
   FA_X1 i_1458 (.A(n_1604), .B(n_1602), .CI(n_1600), .CO(n_1617), .S(n_1616));
   FA_X1 i_1459 (.A(n_1506), .B(n_1504), .CI(n_1502), .CO(n_1619), .S(n_1618));
   FA_X1 i_1460 (.A(n_1606), .B(n_1512), .CI(n_1510), .CO(n_1621), .S(n_1620));
   FA_X1 i_1461 (.A(n_1508), .B(n_1614), .CI(n_1612), .CO(n_1623), .S(n_1622));
   FA_X1 i_1462 (.A(n_1610), .B(n_1608), .CI(n_1514), .CO(n_1625), .S(n_1624));
   FA_X1 i_1463 (.A(n_1618), .B(n_1616), .CI(n_1516), .CO(n_1627), .S(n_1626));
   FA_X1 i_1464 (.A(n_1518), .B(n_1620), .CI(n_1520), .CO(n_1629), .S(n_1628));
   FA_X1 i_1465 (.A(n_1624), .B(n_1622), .CI(n_1522), .CO(n_1631), .S(n_1630));
   FA_X1 i_1466 (.A(n_1626), .B(n_1524), .CI(n_1628), .CO(n_1633), .S(n_1632));
   FA_X1 i_1467 (.A(n_1630), .B(n_1526), .CI(n_1632), .CO(n_1635), .S(n_1634));
   FA_X1 i_1532 (.A(n_1588), .B(n_1581), .CI(n_1574), .CO(n_1701), .S(n_1700));
   FA_X1 i_1533 (.A(n_1567), .B(n_1560), .CI(n_1553), .CO(n_1703), .S(n_1702));
   FA_X1 i_1534 (.A(n_1546), .B(n_1539), .CI(n_1532), .CO(n_1705), .S(n_1704));
   FA_X1 i_1535 (.A(n_1605), .B(n_1603), .CI(n_1601), .CO(n_1707), .S(n_1706));
   FA_X1 i_1536 (.A(n_1595), .B(n_1693), .CI(n_1687), .CO(n_1709), .S(n_1708));
   FA_X1 i_1537 (.A(n_1680), .B(n_1673), .CI(n_1666), .CO(n_1711), .S(n_1710));
   FA_X1 i_1538 (.A(n_1659), .B(n_1652), .CI(n_1645), .CO(n_1713), .S(n_1712));
   FA_X1 i_1539 (.A(n_1638), .B(n_1607), .CI(n_1704), .CO(n_1715), .S(n_1714));
   FA_X1 i_1540 (.A(n_1702), .B(n_1700), .CI(n_1613), .CO(n_1717), .S(n_1716));
   FA_X1 i_1541 (.A(n_1611), .B(n_1609), .CI(n_1615), .CO(n_1719), .S(n_1718));
   FA_X1 i_1542 (.A(n_1706), .B(n_1619), .CI(n_1617), .CO(n_1721), .S(n_1720));
   FA_X1 i_1543 (.A(n_1712), .B(n_1710), .CI(n_1708), .CO(n_1723), .S(n_1722));
   FA_X1 i_1544 (.A(n_1714), .B(n_1621), .CI(n_1718), .CO(n_1725), .S(n_1724));
   FA_X1 i_1545 (.A(n_1716), .B(n_1623), .CI(n_1625), .CO(n_1727), .S(n_1726));
   FA_X1 i_1546 (.A(n_1720), .B(n_1627), .CI(n_1722), .CO(n_1729), .S(n_1728));
   FA_X1 i_1547 (.A(n_1724), .B(n_1629), .CI(n_1726), .CO(n_1731), .S(n_1730));
   FA_X1 i_1548 (.A(n_1631), .B(n_1728), .CI(n_1730), .CO(n_1733), .S(n_1732));
   HA_X1 i_1549 (.A(n_1633), .B(n_1732), .CO(n_1735), .S(n_1734));
   FA_X1 i_1606 (.A(\sums[0] [19]), .B(n_1694), .CI(n_1688), .CO(n_1), .S(n_0));
   FA_X1 i_1607 (.A(n_1681), .B(n_1674), .CI(n_1667), .CO(n_3), .S(n_2));
   FA_X1 i_1608 (.A(n_1660), .B(n_1653), .CI(n_1646), .CO(n_5), .S(n_4));
   FA_X1 i_1609 (.A(n_1639), .B(n_1705), .CI(n_1703), .CO(n_7), .S(n_6));
   FA_X1 i_1610 (.A(n_1701), .B(n_281), .CI(n_280), .CO(n_9), .S(n_8));
   FA_X1 i_1611 (.A(n_1773), .B(n_1766), .CI(n_1759), .CO(n_11), .S(n_10));
   FA_X1 i_1612 (.A(n_1752), .B(n_1745), .CI(n_1738), .CO(n_13), .S(n_12));
   FA_X1 i_1613 (.A(n_1707), .B(n_4), .CI(n_2), .CO(n_15), .S(n_14));
   FA_X1 i_1614 (.A(n_0), .B(n_1713), .CI(n_1711), .CO(n_17), .S(n_16));
   FA_X1 i_1615 (.A(n_1709), .B(n_6), .CI(n_1717), .CO(n_19), .S(n_18));
   FA_X1 i_1616 (.A(n_1715), .B(n_1719), .CI(n_12), .CO(n_21), .S(n_20));
   FA_X1 i_1617 (.A(n_10), .B(n_8), .CI(n_1721), .CO(n_23), .S(n_22));
   FA_X1 i_1618 (.A(n_16), .B(n_14), .CI(n_1723), .CO(n_25), .S(n_24));
   FA_X1 i_1619 (.A(n_18), .B(n_1725), .CI(n_20), .CO(n_27), .S(n_26));
   FA_X1 i_1620 (.A(n_1727), .B(n_22), .CI(n_24), .CO(n_29), .S(n_28));
   FA_X1 i_1621 (.A(n_1729), .B(n_26), .CI(n_1731), .CO(n_31), .S(n_30));
   FA_X1 i_1622 (.A(n_28), .B(n_1733), .CI(n_30), .CO(n_33), .S(n_32));
   FA_X1 i_1680 (.A(n_279), .B(n_1774), .CI(n_1767), .CO(n_35), .S(n_34));
   FA_X1 i_1681 (.A(n_1760), .B(n_1753), .CI(n_1746), .CO(n_37), .S(n_36));
   FA_X1 i_1682 (.A(n_1739), .B(n_5), .CI(n_3), .CO(n_39), .S(n_38));
   FA_X1 i_1683 (.A(n_1), .B(n_278), .CI(n_277), .CO(n_41), .S(n_40));
   FA_X1 i_1684 (.A(n_276), .B(n_275), .CI(n_274), .CO(n_43), .S(n_42));
   FA_X1 i_1685 (.A(n_273), .B(n_272), .CI(n_271), .CO(n_45), .S(n_44));
   FA_X1 i_1686 (.A(n_7), .B(n_36), .CI(n_34), .CO(n_47), .S(n_46));
   FA_X1 i_1687 (.A(n_13), .B(n_11), .CI(n_9), .CO(n_49), .S(n_48));
   FA_X1 i_1688 (.A(n_38), .B(n_17), .CI(n_15), .CO(n_51), .S(n_50));
   FA_X1 i_1689 (.A(n_44), .B(n_42), .CI(n_40), .CO(n_53), .S(n_52));
   FA_X1 i_1690 (.A(n_19), .B(n_48), .CI(n_46), .CO(n_55), .S(n_54));
   FA_X1 i_1691 (.A(n_21), .B(n_23), .CI(n_50), .CO(n_57), .S(n_56));
   FA_X1 i_1692 (.A(n_25), .B(n_52), .CI(n_27), .CO(n_59), .S(n_58));
   FA_X1 i_1693 (.A(n_54), .B(n_56), .CI(n_29), .CO(n_61), .S(n_60));
   FA_X1 i_1694 (.A(n_58), .B(n_31), .CI(n_60), .CO(n_63), .S(n_62));
   FA_X1 i_1745 (.A(n_270), .B(n_269), .CI(n_268), .CO(n_65), .S(n_64));
   FA_X1 i_1746 (.A(n_267), .B(n_266), .CI(n_265), .CO(n_67), .S(n_66));
   FA_X1 i_1747 (.A(n_264), .B(n_37), .CI(n_35), .CO(n_69), .S(n_68));
   FA_X1 i_1748 (.A(n_263), .B(n_261), .CI(n_260), .CO(n_71), .S(n_70));
   FA_X1 i_1749 (.A(n_259), .B(n_258), .CI(n_257), .CO(n_73), .S(n_72));
   FA_X1 i_1750 (.A(n_256), .B(n_255), .CI(n_39), .CO(n_75), .S(n_74));
   FA_X1 i_1751 (.A(n_66), .B(n_64), .CI(n_45), .CO(n_77), .S(n_76));
   FA_X1 i_1752 (.A(n_43), .B(n_41), .CI(n_68), .CO(n_79), .S(n_78));
   FA_X1 i_1753 (.A(n_49), .B(n_47), .CI(n_74), .CO(n_81), .S(n_80));
   FA_X1 i_1754 (.A(n_72), .B(n_70), .CI(n_51), .CO(n_83), .S(n_82));
   FA_X1 i_1755 (.A(n_78), .B(n_76), .CI(n_53), .CO(n_85), .S(n_84));
   FA_X1 i_1756 (.A(n_80), .B(n_55), .CI(n_82), .CO(n_87), .S(n_86));
   FA_X1 i_1757 (.A(n_57), .B(n_84), .CI(n_59), .CO(n_89), .S(n_88));
   FA_X1 i_1758 (.A(n_86), .B(n_61), .CI(n_88), .CO(n_91), .S(n_90));
   FA_X1 i_1801 (.A(\sums[0] [22]), .B(n_262), .CI(n_254), .CO(n_93), .S(n_92));
   FA_X1 i_1802 (.A(n_253), .B(n_252), .CI(n_251), .CO(n_95), .S(n_94));
   FA_X1 i_1803 (.A(n_250), .B(n_249), .CI(n_67), .CO(n_97), .S(n_96));
   FA_X1 i_1804 (.A(n_65), .B(n_248), .CI(n_247), .CO(n_99), .S(n_98));
   FA_X1 i_1805 (.A(n_246), .B(n_245), .CI(n_244), .CO(n_101), .S(n_100));
   FA_X1 i_1806 (.A(n_243), .B(n_69), .CI(n_96), .CO(n_103), .S(n_102));
   FA_X1 i_1807 (.A(n_94), .B(n_92), .CI(n_73), .CO(n_105), .S(n_104));
   FA_X1 i_1808 (.A(n_71), .B(n_75), .CI(n_77), .CO(n_107), .S(n_106));
   FA_X1 i_1809 (.A(n_100), .B(n_98), .CI(n_102), .CO(n_109), .S(n_108));
   FA_X1 i_1810 (.A(n_79), .B(n_104), .CI(n_81), .CO(n_111), .S(n_110));
   FA_X1 i_1811 (.A(n_106), .B(n_83), .CI(n_85), .CO(n_113), .S(n_112));
   FA_X1 i_1812 (.A(n_108), .B(n_110), .CI(n_87), .CO(n_115), .S(n_114));
   FA_X1 i_1813 (.A(n_112), .B(n_89), .CI(n_114), .CO(n_117), .S(n_116));
   FA_X1 i_1857 (.A(n_242), .B(n_241), .CI(n_240), .CO(n_119), .S(n_118));
   FA_X1 i_1858 (.A(n_239), .B(n_238), .CI(n_95), .CO(n_121), .S(n_120));
   FA_X1 i_1859 (.A(n_93), .B(n_237), .CI(n_236), .CO(n_123), .S(n_122));
   FA_X1 i_1860 (.A(n_235), .B(n_234), .CI(n_233), .CO(n_125), .S(n_124));
   FA_X1 i_1861 (.A(n_232), .B(n_97), .CI(n_120), .CO(n_127), .S(n_126));
   FA_X1 i_1862 (.A(n_118), .B(n_101), .CI(n_99), .CO(n_129), .S(n_128));
   FA_X1 i_1863 (.A(n_105), .B(n_103), .CI(n_124), .CO(n_131), .S(n_130));
   FA_X1 i_1864 (.A(n_122), .B(n_126), .CI(n_107), .CO(n_133), .S(n_132));
   FA_X1 i_1865 (.A(n_128), .B(n_109), .CI(n_130), .CO(n_135), .S(n_134));
   FA_X1 i_1866 (.A(n_111), .B(n_132), .CI(n_113), .CO(n_137), .S(n_136));
   FA_X1 i_1867 (.A(n_134), .B(n_115), .CI(n_136), .CO(n_139), .S(n_138));
   FA_X1 i_1904 (.A(n_231), .B(n_230), .CI(n_229), .CO(n_141), .S(n_140));
   FA_X1 i_1905 (.A(n_228), .B(n_227), .CI(n_119), .CO(n_143), .S(n_142));
   FA_X1 i_1906 (.A(n_226), .B(n_224), .CI(n_223), .CO(n_145), .S(n_144));
   FA_X1 i_1907 (.A(n_222), .B(n_221), .CI(n_220), .CO(n_147), .S(n_146));
   FA_X1 i_1908 (.A(n_121), .B(n_142), .CI(n_140), .CO(n_149), .S(n_148));
   FA_X1 i_1909 (.A(n_125), .B(n_123), .CI(n_129), .CO(n_151), .S(n_150));
   FA_X1 i_1910 (.A(n_127), .B(n_146), .CI(n_144), .CO(n_153), .S(n_152));
   FA_X1 i_1911 (.A(n_150), .B(n_148), .CI(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_1912 (.A(n_133), .B(n_152), .CI(n_135), .CO(n_157), .S(n_156));
   FA_X1 i_1913 (.A(n_154), .B(n_137), .CI(n_156), .CO(n_159), .S(n_158));
   FA_X1 i_1942 (.A(\sums[0] [25]), .B(n_225), .CI(n_219), .CO(n_161), .S(n_160));
   FA_X1 i_1943 (.A(n_218), .B(n_217), .CI(n_216), .CO(n_163), .S(n_162));
   FA_X1 i_1944 (.A(n_141), .B(n_215), .CI(n_214), .CO(n_165), .S(n_164));
   FA_X1 i_1945 (.A(n_213), .B(n_212), .CI(n_143), .CO(n_167), .S(n_166));
   FA_X1 i_1946 (.A(n_162), .B(n_160), .CI(n_147), .CO(n_169), .S(n_168));
   FA_X1 i_1947 (.A(n_145), .B(n_149), .CI(n_166), .CO(n_171), .S(n_170));
   FA_X1 i_1948 (.A(n_164), .B(n_151), .CI(n_168), .CO(n_173), .S(n_172));
   FA_X1 i_1949 (.A(n_153), .B(n_170), .CI(n_155), .CO(n_175), .S(n_174));
   FA_X1 i_1950 (.A(n_172), .B(n_157), .CI(n_174), .CO(n_177), .S(n_176));
   FA_X1 i_1983 (.A(n_501), .B(n_513), .CI(n_211), .CO(n_179), .S(n_178));
   FA_X1 i_1984 (.A(n_539), .B(n_537), .CI(n_179), .CO(n_181), .S(n_180));
   FA_X1 i_1985 (.A(n_572), .B(n_574), .CI(n_181), .CO(n_183), .S(n_182));
   FA_X1 i_1986 (.A(n_612), .B(n_610), .CI(n_183), .CO(n_185), .S(n_184));
   FA_X1 i_1987 (.A(n_660), .B(n_658), .CI(n_185), .CO(n_187), .S(n_186));
   FA_X1 i_1988 (.A(n_715), .B(n_717), .CI(n_187), .CO(n_189), .S(n_188));
   FA_X1 i_1989 (.A(n_775), .B(n_777), .CI(n_189), .CO(n_191), .S(n_190));
   FA_X1 i_1990 (.A(n_847), .B(n_845), .CI(n_191), .CO(n_193), .S(n_192));
   FA_X1 i_1991 (.A(n_924), .B(n_926), .CI(n_193), .CO(n_195), .S(n_194));
   FA_X1 i_1992 (.A(n_1006), .B(n_1008), .CI(n_195), .CO(n_196), .S(
      \sums[2] [11]));
   FA_X1 i_1993 (.A(n_1009), .B(n_1100), .CI(n_196), .CO(n_197), .S(
      \sums[2] [12]));
   FA_X1 i_1994 (.A(n_1101), .B(n_1201), .CI(n_197), .CO(n_198), .S(
      \sums[2] [13]));
   FA_X1 i_1995 (.A(n_1202), .B(n_1305), .CI(n_198), .CO(n_199), .S(
      \sums[2] [14]));
   FA_X1 i_1996 (.A(n_1306), .B(n_1419), .CI(n_199), .CO(n_200), .S(
      \sums[2] [15]));
   FA_X1 i_1997 (.A(n_1420), .B(n_1527), .CI(n_200), .CO(n_201), .S(
      \sums[2] [16]));
   FA_X1 i_1998 (.A(n_1528), .B(n_1634), .CI(n_201), .CO(n_202), .S(
      \sums[2] [17]));
   FA_X1 i_1999 (.A(n_1635), .B(n_1734), .CI(n_202), .CO(n_203), .S(
      \sums[2] [18]));
   FA_X1 i_2000 (.A(n_1735), .B(n_32), .CI(n_203), .CO(n_204), .S(\sums[2] [19]));
   FA_X1 i_2001 (.A(n_62), .B(n_33), .CI(n_204), .CO(n_205), .S(\sums[2] [20]));
   FA_X1 i_2002 (.A(n_63), .B(n_90), .CI(n_205), .CO(n_206), .S(\sums[2] [21]));
   FA_X1 i_2003 (.A(n_91), .B(n_116), .CI(n_206), .CO(n_207), .S(\sums[2] [22]));
   FA_X1 i_2004 (.A(n_138), .B(n_117), .CI(n_207), .CO(n_208), .S(\sums[2] [23]));
   FA_X1 i_2005 (.A(n_139), .B(n_158), .CI(n_208), .CO(n_209), .S(\sums[2] [24]));
   FA_X1 i_2006 (.A(n_159), .B(n_176), .CI(n_209), .CO(n_210), .S(\sums[2] [25]));
   NOR2_X1 i_0 (.A1(n_284), .A2(n_282), .ZN(n_211));
   AOI21_X1 i_1 (.A(n_283), .B1(\r_weights[1] [1]), .B2(n_285), .ZN(n_282));
   XOR2_X1 i_2 (.A(n_1648), .B(n_1647), .Z(n_283));
   AOI21_X1 i_3 (.A(n_285), .B1(\r_values[1] [0]), .B2(\r_weights[1] [1]), 
      .ZN(n_284));
   AND4_X1 i_4 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [0]), .A3(
      \r_values[1] [0]), .A4(\r_weights[1] [0]), .ZN(n_285));
   XOR2_X1 i_5 (.A(n_1593), .B(n_286), .Z(n_501));
   NAND2_X1 i_6 (.A1(n_1597), .A2(n_1596), .ZN(n_286));
   XOR2_X1 i_7 (.A(n_1668), .B(n_287), .Z(n_212));
   NAND2_X1 i_8 (.A1(n_1671), .A2(n_1669), .ZN(n_287));
   XOR2_X1 i_9 (.A(n_1677), .B(n_288), .Z(n_213));
   NAND2_X1 i_10 (.A1(n_1682), .A2(n_1678), .ZN(n_288));
   XNOR2_X1 i_11 (.A(n_1656), .B(n_289), .ZN(n_214));
   NAND2_X1 i_12 (.A1(n_1662), .A2(n_1658), .ZN(n_289));
   XNOR2_X1 i_13 (.A(n_1685), .B(n_290), .ZN(n_215));
   NAND2_X1 i_14 (.A1(n_1691), .A2(n_1689), .ZN(n_290));
   OAI21_X1 i_15 (.A(n_292), .B1(n_295), .B2(n_294), .ZN(n_216));
   OAI21_X1 i_16 (.A(n_297), .B1(n_300), .B2(n_299), .ZN(n_217));
   AOI21_X1 i_17 (.A(n_303), .B1(n_305), .B2(n_304), .ZN(n_218));
   OAI22_X1 i_18 (.A1(n_1686), .A2(n_357), .B1(n_1664), .B2(n_307), .ZN(n_219));
   XOR2_X1 i_19 (.A(n_295), .B(n_291), .Z(n_220));
   NAND2_X1 i_20 (.A1(n_293), .A2(n_292), .ZN(n_291));
   NAND3_X1 i_21 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [10]), .A3(n_1672), 
      .ZN(n_292));
   INV_X1 i_22 (.A(n_294), .ZN(n_293));
   AOI21_X1 i_23 (.A(n_1672), .B1(\r_values[0] [14]), .B2(\r_weights[0] [10]), 
      .ZN(n_294));
   NAND2_X1 i_24 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [9]), .ZN(n_295));
   XOR2_X1 i_25 (.A(n_300), .B(n_296), .Z(n_221));
   NAND2_X1 i_26 (.A1(n_298), .A2(n_297), .ZN(n_296));
   NAND3_X1 i_27 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [13]), .A3(n_1683), 
      .ZN(n_297));
   INV_X1 i_28 (.A(n_299), .ZN(n_298));
   AOI21_X1 i_29 (.A(n_1683), .B1(\r_values[0] [11]), .B2(\r_weights[0] [13]), 
      .ZN(n_299));
   NAND2_X1 i_30 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [12]), .ZN(n_300));
   XOR2_X1 i_31 (.A(n_305), .B(n_301), .Z(n_222));
   NAND2_X1 i_32 (.A1(n_304), .A2(n_302), .ZN(n_301));
   INV_X1 i_33 (.A(n_303), .ZN(n_302));
   AOI22_X1 i_34 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [10]), .B1(
      \r_values[1] [15]), .B2(\r_weights[1] [9]), .ZN(n_303));
   NAND2_X1 i_35 (.A1(n_1656), .A2(n_352), .ZN(n_304));
   NAND2_X1 i_36 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [15]), .ZN(n_305));
   XOR2_X1 i_37 (.A(n_1663), .B(n_306), .Z(n_223));
   AOI21_X1 i_38 (.A(n_307), .B1(n_1685), .B2(n_356), .ZN(n_306));
   AOI22_X1 i_39 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [13]), .B1(
      \r_values[1] [12]), .B2(\r_weights[1] [12]), .ZN(n_307));
   OAI21_X1 i_40 (.A(n_308), .B1(n_311), .B2(n_225), .ZN(n_224));
   OAI21_X1 i_41 (.A(\sums[0] [24]), .B1(n_311), .B2(n_309), .ZN(n_308));
   OAI21_X1 i_42 (.A(n_310), .B1(n_1778), .B2(n_311), .ZN(n_225));
   INV_X1 i_43 (.A(n_310), .ZN(n_309));
   NAND3_X1 i_44 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [15]), .A3(n_1692), 
      .ZN(n_310));
   AOI21_X1 i_45 (.A(n_1692), .B1(\r_values[1] [9]), .B2(\r_weights[1] [15]), 
      .ZN(n_311));
   INV_X1 i_46 (.A(n_312), .ZN(n_226));
   AOI22_X1 i_47 (.A1(\sums[0] [23]), .A2(n_362), .B1(n_334), .B2(n_333), 
      .ZN(n_312));
   OAI21_X1 i_48 (.A(n_314), .B1(n_317), .B2(n_316), .ZN(n_227));
   OAI21_X1 i_49 (.A(n_319), .B1(n_322), .B2(n_321), .ZN(n_228));
   AOI21_X1 i_50 (.A(n_326), .B1(n_327), .B2(n_324), .ZN(n_229));
   OAI22_X1 i_51 (.A1(n_1664), .A2(n_389), .B1(n_353), .B2(n_329), .ZN(n_230));
   OAI21_X1 i_52 (.A(n_331), .B1(n_357), .B2(n_332), .ZN(n_231));
   XOR2_X1 i_53 (.A(n_317), .B(n_313), .Z(n_232));
   NAND2_X1 i_54 (.A1(n_315), .A2(n_314), .ZN(n_313));
   NAND4_X1 i_55 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [9]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [10]), .ZN(n_314));
   INV_X1 i_56 (.A(n_316), .ZN(n_315));
   AOI22_X1 i_57 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [9]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [10]), .ZN(n_316));
   NAND2_X1 i_58 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [8]), .ZN(n_317));
   XOR2_X1 i_59 (.A(n_322), .B(n_318), .Z(n_233));
   NAND2_X1 i_60 (.A1(n_320), .A2(n_319), .ZN(n_318));
   NAND4_X1 i_61 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [12]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [13]), .ZN(n_319));
   INV_X1 i_62 (.A(n_321), .ZN(n_320));
   AOI22_X1 i_63 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [12]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [13]), .ZN(n_321));
   NAND2_X1 i_64 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [11]), .ZN(n_322));
   XOR2_X1 i_65 (.A(n_327), .B(n_323), .Z(n_234));
   NAND2_X1 i_66 (.A1(n_325), .A2(n_324), .ZN(n_323));
   NAND3_X1 i_67 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [8]), .A3(n_347), 
      .ZN(n_324));
   INV_X1 i_68 (.A(n_326), .ZN(n_325));
   AOI21_X1 i_69 (.A(n_347), .B1(\r_values[1] [15]), .B2(\r_weights[1] [8]), 
      .ZN(n_326));
   NAND2_X1 i_70 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [14]), .ZN(n_327));
   XOR2_X1 i_71 (.A(n_352), .B(n_328), .Z(n_235));
   AOI21_X1 i_72 (.A(n_329), .B1(n_1663), .B2(n_388), .ZN(n_328));
   AOI22_X1 i_73 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [11]), .B1(
      \r_values[1] [13]), .B2(\r_weights[1] [10]), .ZN(n_329));
   XOR2_X1 i_74 (.A(n_356), .B(n_330), .Z(n_236));
   AOI21_X1 i_75 (.A(n_332), .B1(n_1692), .B2(n_392), .ZN(n_330));
   NAND2_X1 i_76 (.A1(n_1692), .A2(n_392), .ZN(n_331));
   AOI22_X1 i_77 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [14]), .B1(
      \r_values[1] [10]), .B2(\r_weights[1] [13]), .ZN(n_332));
   XOR2_X1 i_78 (.A(n_334), .B(n_333), .Z(n_237));
   OAI21_X1 i_79 (.A(n_361), .B1(n_393), .B2(n_360), .ZN(n_333));
   XNOR2_X1 i_80 (.A(\sums[0] [23]), .B(n_363), .ZN(n_334));
   OAI21_X1 i_81 (.A(n_336), .B1(n_339), .B2(n_338), .ZN(n_238));
   OAI21_X1 i_82 (.A(n_341), .B1(n_344), .B2(n_343), .ZN(n_239));
   OAI21_X1 i_83 (.A(n_346), .B1(n_350), .B2(n_349), .ZN(n_240));
   OAI22_X1 i_84 (.A1(n_422), .A2(n_353), .B1(n_385), .B2(n_354), .ZN(n_241));
   OAI22_X1 i_85 (.A1(n_426), .A2(n_357), .B1(n_389), .B2(n_358), .ZN(n_242));
   XOR2_X1 i_86 (.A(n_339), .B(n_335), .Z(n_243));
   NAND2_X1 i_87 (.A1(n_337), .A2(n_336), .ZN(n_335));
   NAND4_X1 i_88 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [8]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [9]), .ZN(n_336));
   INV_X1 i_89 (.A(n_338), .ZN(n_337));
   AOI22_X1 i_90 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [9]), .ZN(n_338));
   NAND2_X1 i_91 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [7]), .ZN(n_339));
   XOR2_X1 i_92 (.A(n_344), .B(n_340), .Z(n_244));
   NAND2_X1 i_93 (.A1(n_342), .A2(n_341), .ZN(n_340));
   NAND4_X1 i_94 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [11]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [12]), .ZN(n_341));
   INV_X1 i_95 (.A(n_343), .ZN(n_342));
   AOI22_X1 i_96 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [11]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [12]), .ZN(n_343));
   NAND2_X1 i_97 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [10]), .ZN(n_344));
   XOR2_X1 i_98 (.A(n_350), .B(n_345), .Z(n_245));
   NAND2_X1 i_99 (.A1(n_348), .A2(n_346), .ZN(n_345));
   NAND2_X1 i_100 (.A1(n_378), .A2(n_347), .ZN(n_346));
   AND2_X1 i_101 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [15]), .ZN(n_347));
   INV_X1 i_102 (.A(n_349), .ZN(n_348));
   AOI22_X1 i_103 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [14]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [15]), .ZN(n_349));
   NAND2_X1 i_104 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [13]), .ZN(n_350));
   XOR2_X1 i_105 (.A(n_384), .B(n_351), .Z(n_246));
   AOI21_X1 i_106 (.A(n_354), .B1(n_421), .B2(n_352), .ZN(n_351));
   INV_X1 i_107 (.A(n_353), .ZN(n_352));
   NAND2_X1 i_108 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [9]), .ZN(n_353));
   AOI22_X1 i_109 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [9]), .B1(
      \r_values[1] [14]), .B2(\r_weights[1] [8]), .ZN(n_354));
   XOR2_X1 i_110 (.A(n_388), .B(n_355), .Z(n_247));
   AOI21_X1 i_111 (.A(n_358), .B1(n_425), .B2(n_356), .ZN(n_355));
   INV_X1 i_112 (.A(n_357), .ZN(n_356));
   NAND2_X1 i_113 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [12]), .ZN(n_357));
   AOI22_X1 i_114 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [12]), .B1(
      \r_values[1] [11]), .B2(\r_weights[1] [11]), .ZN(n_358));
   XOR2_X1 i_115 (.A(n_392), .B(n_359), .Z(n_248));
   AOI21_X1 i_116 (.A(n_360), .B1(n_430), .B2(n_362), .ZN(n_359));
   AOI22_X1 i_117 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [15]), .B1(
      \r_values[1] [8]), .B2(\r_weights[1] [14]), .ZN(n_360));
   NAND2_X1 i_118 (.A1(n_430), .A2(n_362), .ZN(n_361));
   INV_X1 i_119 (.A(n_363), .ZN(n_362));
   NAND2_X1 i_120 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [15]), .ZN(n_363));
   OAI21_X1 i_121 (.A(n_365), .B1(n_368), .B2(n_367), .ZN(n_249));
   OAI21_X1 i_122 (.A(n_370), .B1(n_373), .B2(n_372), .ZN(n_250));
   OAI21_X1 i_123 (.A(n_375), .B1(n_379), .B2(n_377), .ZN(n_251));
   AOI21_X1 i_124 (.A(n_382), .B1(n_386), .B2(n_383), .ZN(n_252));
   OAI22_X1 i_125 (.A1(n_461), .A2(n_389), .B1(n_422), .B2(n_390), .ZN(n_253));
   OAI22_X1 i_126 (.A1(n_465), .A2(n_393), .B1(n_426), .B2(n_394), .ZN(n_254));
   XOR2_X1 i_127 (.A(n_368), .B(n_364), .Z(n_255));
   NAND2_X1 i_128 (.A1(n_366), .A2(n_365), .ZN(n_364));
   NAND4_X1 i_129 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [7]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [8]), .ZN(n_365));
   INV_X1 i_130 (.A(n_367), .ZN(n_366));
   AOI22_X1 i_131 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [7]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [8]), .ZN(n_367));
   NAND2_X1 i_132 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [6]), .ZN(n_368));
   XOR2_X1 i_133 (.A(n_373), .B(n_369), .Z(n_256));
   NAND2_X1 i_134 (.A1(n_371), .A2(n_370), .ZN(n_369));
   NAND4_X1 i_135 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [10]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [11]), .ZN(n_370));
   INV_X1 i_136 (.A(n_372), .ZN(n_371));
   AOI22_X1 i_137 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [10]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [11]), .ZN(n_372));
   NAND2_X1 i_138 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [9]), .ZN(n_373));
   XOR2_X1 i_139 (.A(n_379), .B(n_374), .Z(n_257));
   NAND2_X1 i_140 (.A1(n_376), .A2(n_375), .ZN(n_374));
   NAND3_X1 i_141 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [13]), .A3(n_378), 
      .ZN(n_375));
   INV_X1 i_142 (.A(n_377), .ZN(n_376));
   AOI21_X1 i_143 (.A(n_378), .B1(\r_values[0] [8]), .B2(\r_weights[0] [13]), 
      .ZN(n_377));
   AND2_X1 i_144 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [14]), .ZN(n_378));
   NAND2_X1 i_145 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [12]), .ZN(n_379));
   XOR2_X1 i_146 (.A(n_386), .B(n_380), .Z(n_258));
   NAND2_X1 i_147 (.A1(n_383), .A2(n_381), .ZN(n_380));
   INV_X1 i_148 (.A(n_382), .ZN(n_381));
   AOI22_X1 i_149 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [7]), .B1(
      \r_values[1] [15]), .B2(\r_weights[1] [6]), .ZN(n_382));
   NAND2_X1 i_150 (.A1(n_456), .A2(n_384), .ZN(n_383));
   INV_X1 i_151 (.A(n_385), .ZN(n_384));
   NAND2_X1 i_152 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [7]), .ZN(n_385));
   NAND2_X1 i_153 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [15]), .ZN(n_386));
   XOR2_X1 i_154 (.A(n_421), .B(n_387), .Z(n_259));
   AOI21_X1 i_155 (.A(n_390), .B1(n_460), .B2(n_388), .ZN(n_387));
   INV_X1 i_156 (.A(n_389), .ZN(n_388));
   NAND2_X1 i_157 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [10]), .ZN(n_389));
   AOI22_X1 i_158 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [10]), .B1(
      \r_values[1] [12]), .B2(\r_weights[1] [9]), .ZN(n_390));
   XOR2_X1 i_159 (.A(n_425), .B(n_391), .Z(n_260));
   AOI21_X1 i_160 (.A(n_394), .B1(n_464), .B2(n_392), .ZN(n_391));
   INV_X1 i_161 (.A(n_393), .ZN(n_392));
   NAND2_X1 i_162 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [13]), .ZN(n_393));
   AOI22_X1 i_163 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [13]), .B1(
      \r_values[1] [9]), .B2(\r_weights[1] [12]), .ZN(n_394));
   AOI21_X1 i_164 (.A(n_395), .B1(n_397), .B2(n_262), .ZN(n_261));
   INV_X1 i_165 (.A(n_396), .ZN(n_395));
   OAI21_X1 i_166 (.A(n_1777), .B1(n_398), .B2(n_262), .ZN(n_396));
   AOI21_X1 i_167 (.A(n_398), .B1(n_1777), .B2(n_397), .ZN(n_262));
   NAND3_X1 i_168 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [15]), .A3(n_430), 
      .ZN(n_397));
   AOI21_X1 i_169 (.A(n_430), .B1(\r_values[1] [6]), .B2(\r_weights[1] [15]), 
      .ZN(n_398));
   INV_X1 i_170 (.A(n_399), .ZN(n_263));
   AOI22_X1 i_171 (.A1(\sums[0] [20]), .A2(n_470), .B1(n_433), .B2(n_432), 
      .ZN(n_399));
   OAI21_X1 i_172 (.A(n_401), .B1(n_404), .B2(n_403), .ZN(n_264));
   OAI21_X1 i_173 (.A(n_406), .B1(n_409), .B2(n_408), .ZN(n_265));
   OAI21_X1 i_174 (.A(n_411), .B1(n_414), .B2(n_413), .ZN(n_266));
   AOI21_X1 i_175 (.A(n_418), .B1(n_419), .B2(n_416), .ZN(n_267));
   OAI22_X1 i_176 (.A1(n_505), .A2(n_422), .B1(n_457), .B2(n_423), .ZN(n_268));
   OAI22_X1 i_177 (.A1(n_510), .A2(n_426), .B1(n_461), .B2(n_427), .ZN(n_269));
   OAI21_X1 i_178 (.A(n_429), .B1(n_465), .B2(n_431), .ZN(n_270));
   XOR2_X1 i_179 (.A(n_404), .B(n_400), .Z(n_271));
   NAND2_X1 i_180 (.A1(n_402), .A2(n_401), .ZN(n_400));
   NAND4_X1 i_181 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [6]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [7]), .ZN(n_401));
   INV_X1 i_182 (.A(n_403), .ZN(n_402));
   AOI22_X1 i_183 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [6]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [7]), .ZN(n_403));
   NAND2_X1 i_184 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [5]), .ZN(n_404));
   XOR2_X1 i_185 (.A(n_409), .B(n_405), .Z(n_272));
   NAND2_X1 i_186 (.A1(n_407), .A2(n_406), .ZN(n_405));
   NAND4_X1 i_187 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [9]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [10]), .ZN(n_406));
   INV_X1 i_188 (.A(n_408), .ZN(n_407));
   AOI22_X1 i_189 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [9]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [10]), .ZN(n_408));
   NAND2_X1 i_190 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [8]), .ZN(n_409));
   XOR2_X1 i_191 (.A(n_414), .B(n_410), .Z(n_273));
   NAND2_X1 i_192 (.A1(n_412), .A2(n_411), .ZN(n_410));
   NAND4_X1 i_193 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [12]), .A3(
      \r_values[0] [7]), .A4(\r_weights[0] [13]), .ZN(n_411));
   INV_X1 i_194 (.A(n_413), .ZN(n_412));
   AOI22_X1 i_195 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [12]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [13]), .ZN(n_413));
   NAND2_X1 i_196 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [11]), .ZN(n_414));
   XOR2_X1 i_197 (.A(n_419), .B(n_415), .Z(n_274));
   NAND2_X1 i_198 (.A1(n_417), .A2(n_416), .ZN(n_415));
   NAND3_X1 i_199 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [5]), .A3(n_451), 
      .ZN(n_416));
   INV_X1 i_200 (.A(n_418), .ZN(n_417));
   AOI21_X1 i_201 (.A(n_451), .B1(\r_values[1] [15]), .B2(\r_weights[1] [5]), 
      .ZN(n_418));
   NAND2_X1 i_202 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [14]), .ZN(n_419));
   XOR2_X1 i_203 (.A(n_456), .B(n_420), .Z(n_275));
   AOI21_X1 i_204 (.A(n_423), .B1(n_504), .B2(n_421), .ZN(n_420));
   INV_X1 i_205 (.A(n_422), .ZN(n_421));
   NAND2_X1 i_206 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [8]), .ZN(n_422));
   AOI22_X1 i_207 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [8]), .B1(
      \r_values[1] [13]), .B2(\r_weights[1] [7]), .ZN(n_423));
   XOR2_X1 i_208 (.A(n_460), .B(n_424), .Z(n_276));
   AOI21_X1 i_209 (.A(n_427), .B1(n_509), .B2(n_425), .ZN(n_424));
   INV_X1 i_210 (.A(n_426), .ZN(n_425));
   NAND2_X1 i_211 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [11]), .ZN(n_426));
   AOI22_X1 i_212 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [11]), .B1(
      \r_values[1] [10]), .B2(\r_weights[1] [10]), .ZN(n_427));
   XOR2_X1 i_213 (.A(n_464), .B(n_428), .Z(n_277));
   AOI21_X1 i_214 (.A(n_431), .B1(n_515), .B2(n_430), .ZN(n_428));
   NAND2_X1 i_215 (.A1(n_515), .A2(n_430), .ZN(n_429));
   AND2_X1 i_216 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [14]), .ZN(n_430));
   AOI22_X1 i_217 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [14]), .B1(
      \r_values[1] [7]), .B2(\r_weights[1] [13]), .ZN(n_431));
   XOR2_X1 i_218 (.A(n_433), .B(n_432), .Z(n_278));
   OAI21_X1 i_219 (.A(n_469), .B1(n_516), .B2(n_468), .ZN(n_432));
   XNOR2_X1 i_220 (.A(\sums[0] [20]), .B(n_471), .ZN(n_433));
   OAI21_X1 i_221 (.A(n_435), .B1(n_438), .B2(n_437), .ZN(n_1739));
   OAI21_X1 i_222 (.A(n_440), .B1(n_443), .B2(n_442), .ZN(n_1746));
   OAI21_X1 i_223 (.A(n_445), .B1(n_448), .B2(n_447), .ZN(n_1753));
   OAI21_X1 i_224 (.A(n_450), .B1(n_454), .B2(n_453), .ZN(n_1760));
   OAI22_X1 i_225 (.A1(n_566), .A2(n_457), .B1(n_499), .B2(n_458), .ZN(n_1767));
   OAI22_X1 i_226 (.A1(n_576), .A2(n_461), .B1(n_505), .B2(n_462), .ZN(n_1774));
   OAI22_X1 i_227 (.A1(n_582), .A2(n_465), .B1(n_510), .B2(n_466), .ZN(n_279));
   XOR2_X1 i_228 (.A(n_438), .B(n_434), .Z(n_1738));
   NAND2_X1 i_229 (.A1(n_436), .A2(n_435), .ZN(n_434));
   NAND4_X1 i_230 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [6]), .ZN(n_435));
   INV_X1 i_231 (.A(n_437), .ZN(n_436));
   AOI22_X1 i_232 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [6]), .ZN(n_437));
   NAND2_X1 i_233 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [4]), .ZN(n_438));
   XOR2_X1 i_234 (.A(n_443), .B(n_439), .Z(n_1745));
   NAND2_X1 i_235 (.A1(n_441), .A2(n_440), .ZN(n_439));
   NAND4_X1 i_236 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [8]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [9]), .ZN(n_440));
   INV_X1 i_237 (.A(n_442), .ZN(n_441));
   AOI22_X1 i_238 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [9]), .ZN(n_442));
   NAND2_X1 i_239 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [7]), .ZN(n_443));
   XOR2_X1 i_240 (.A(n_448), .B(n_444), .Z(n_1752));
   NAND2_X1 i_241 (.A1(n_446), .A2(n_445), .ZN(n_444));
   NAND4_X1 i_242 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [11]), .A3(
      \r_values[0] [7]), .A4(\r_weights[0] [12]), .ZN(n_445));
   INV_X1 i_243 (.A(n_447), .ZN(n_446));
   AOI22_X1 i_244 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [11]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [12]), .ZN(n_447));
   NAND2_X1 i_245 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [10]), .ZN(n_448));
   XOR2_X1 i_246 (.A(n_454), .B(n_449), .Z(n_1759));
   NAND2_X1 i_247 (.A1(n_452), .A2(n_450), .ZN(n_449));
   NAND2_X1 i_248 (.A1(n_491), .A2(n_451), .ZN(n_450));
   AND2_X1 i_249 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [15]), .ZN(n_451));
   INV_X1 i_250 (.A(n_453), .ZN(n_452));
   AOI22_X1 i_251 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [14]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [15]), .ZN(n_453));
   NAND2_X1 i_252 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [13]), .ZN(n_454));
   XOR2_X1 i_253 (.A(n_498), .B(n_455), .Z(n_1766));
   AOI21_X1 i_254 (.A(n_458), .B1(n_563), .B2(n_456), .ZN(n_455));
   INV_X1 i_255 (.A(n_457), .ZN(n_456));
   NAND2_X1 i_256 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [6]), .ZN(n_457));
   AOI22_X1 i_257 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [6]), .B1(
      \r_values[1] [14]), .B2(\r_weights[1] [5]), .ZN(n_458));
   XOR2_X1 i_258 (.A(n_504), .B(n_459), .Z(n_1773));
   AOI21_X1 i_259 (.A(n_462), .B1(n_569), .B2(n_460), .ZN(n_459));
   INV_X1 i_260 (.A(n_461), .ZN(n_460));
   NAND2_X1 i_261 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [9]), .ZN(n_461));
   AOI22_X1 i_262 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [9]), .B1(
      \r_values[1] [11]), .B2(\r_weights[1] [8]), .ZN(n_462));
   XOR2_X1 i_263 (.A(n_509), .B(n_463), .Z(n_280));
   AOI21_X1 i_264 (.A(n_466), .B1(n_581), .B2(n_464), .ZN(n_463));
   INV_X1 i_265 (.A(n_465), .ZN(n_464));
   NAND2_X1 i_266 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [12]), .ZN(n_465));
   AOI22_X1 i_267 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [12]), .B1(
      \r_values[1] [8]), .B2(\r_weights[1] [11]), .ZN(n_466));
   XOR2_X1 i_268 (.A(n_515), .B(n_467), .Z(n_281));
   AOI21_X1 i_269 (.A(n_468), .B1(n_588), .B2(n_470), .ZN(n_467));
   AOI22_X1 i_270 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [15]), .B1(
      \r_values[1] [5]), .B2(\r_weights[1] [14]), .ZN(n_468));
   NAND2_X1 i_271 (.A1(n_588), .A2(n_470), .ZN(n_469));
   INV_X1 i_272 (.A(n_471), .ZN(n_470));
   NAND2_X1 i_273 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [15]), .ZN(n_471));
   OAI21_X1 i_274 (.A(n_473), .B1(n_476), .B2(n_475), .ZN(n_1639));
   OAI21_X1 i_275 (.A(n_478), .B1(n_481), .B2(n_480), .ZN(n_1646));
   OAI21_X1 i_276 (.A(n_483), .B1(n_486), .B2(n_485), .ZN(n_1653));
   OAI21_X1 i_277 (.A(n_488), .B1(n_492), .B2(n_490), .ZN(n_1660));
   AOI21_X1 i_278 (.A(n_496), .B1(n_500), .B2(n_497), .ZN(n_1667));
   OAI22_X1 i_279 (.A1(n_649), .A2(n_505), .B1(n_566), .B2(n_506), .ZN(n_1674));
   OAI22_X1 i_280 (.A1(n_667), .A2(n_510), .B1(n_576), .B2(n_511), .ZN(n_1681));
   OAI22_X1 i_281 (.A1(n_673), .A2(n_516), .B1(n_582), .B2(n_518), .ZN(n_1688));
   XOR2_X1 i_282 (.A(n_476), .B(n_472), .Z(n_1638));
   NAND2_X1 i_283 (.A1(n_474), .A2(n_473), .ZN(n_472));
   NAND4_X1 i_284 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [4]), .A3(
      \r_values[0] [13]), .A4(\r_weights[0] [5]), .ZN(n_473));
   INV_X1 i_285 (.A(n_475), .ZN(n_474));
   AOI22_X1 i_286 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [4]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [5]), .ZN(n_475));
   NAND2_X1 i_287 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [3]), .ZN(n_476));
   XOR2_X1 i_288 (.A(n_481), .B(n_477), .Z(n_1645));
   NAND2_X1 i_289 (.A1(n_479), .A2(n_478), .ZN(n_477));
   NAND4_X1 i_290 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [7]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [8]), .ZN(n_478));
   INV_X1 i_291 (.A(n_480), .ZN(n_479));
   AOI22_X1 i_292 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [7]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [8]), .ZN(n_480));
   NAND2_X1 i_293 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [6]), .ZN(n_481));
   XOR2_X1 i_294 (.A(n_486), .B(n_482), .Z(n_1652));
   NAND2_X1 i_295 (.A1(n_484), .A2(n_483), .ZN(n_482));
   NAND4_X1 i_296 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [10]), .A3(
      \r_values[0] [7]), .A4(\r_weights[0] [11]), .ZN(n_483));
   INV_X1 i_297 (.A(n_485), .ZN(n_484));
   AOI22_X1 i_298 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [10]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [11]), .ZN(n_485));
   NAND2_X1 i_299 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [9]), .ZN(n_486));
   XOR2_X1 i_300 (.A(n_492), .B(n_487), .Z(n_1659));
   NAND2_X1 i_301 (.A1(n_489), .A2(n_488), .ZN(n_487));
   NAND3_X1 i_302 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [13]), .A3(n_491), 
      .ZN(n_488));
   INV_X1 i_303 (.A(n_490), .ZN(n_489));
   AOI21_X1 i_304 (.A(n_491), .B1(\r_values[0] [5]), .B2(\r_weights[0] [13]), 
      .ZN(n_490));
   AND2_X1 i_305 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [14]), .ZN(n_491));
   NAND2_X1 i_306 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [12]), .ZN(n_492));
   XOR2_X1 i_307 (.A(n_500), .B(n_493), .Z(n_1666));
   NAND2_X1 i_308 (.A1(n_497), .A2(n_494), .ZN(n_493));
   INV_X1 i_309 (.A(n_496), .ZN(n_494));
   AOI22_X1 i_310 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [4]), .B1(
      \r_values[1] [15]), .B2(\r_weights[1] [3]), .ZN(n_496));
   NAND2_X1 i_311 (.A1(n_642), .A2(n_498), .ZN(n_497));
   INV_X1 i_312 (.A(n_499), .ZN(n_498));
   NAND2_X1 i_313 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [4]), .ZN(n_499));
   NAND2_X1 i_314 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [15]), .ZN(n_500));
   XOR2_X1 i_315 (.A(n_563), .B(n_503), .Z(n_1673));
   AOI21_X1 i_316 (.A(n_506), .B1(n_648), .B2(n_504), .ZN(n_503));
   INV_X1 i_317 (.A(n_505), .ZN(n_504));
   NAND2_X1 i_318 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [7]), .ZN(n_505));
   AOI22_X1 i_319 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [7]), .B1(
      \r_values[1] [12]), .B2(\r_weights[1] [6]), .ZN(n_506));
   XOR2_X1 i_320 (.A(n_569), .B(n_507), .Z(n_1680));
   AOI21_X1 i_321 (.A(n_511), .B1(n_666), .B2(n_509), .ZN(n_507));
   INV_X1 i_322 (.A(n_510), .ZN(n_509));
   NAND2_X1 i_323 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [10]), .ZN(n_510));
   AOI22_X1 i_324 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [10]), .B1(
      \r_values[1] [9]), .B2(\r_weights[1] [9]), .ZN(n_511));
   XOR2_X1 i_325 (.A(n_581), .B(n_512), .Z(n_1687));
   AOI21_X1 i_326 (.A(n_518), .B1(n_670), .B2(n_515), .ZN(n_512));
   INV_X1 i_327 (.A(n_516), .ZN(n_515));
   NAND2_X1 i_328 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [13]), .ZN(n_516));
   AOI22_X1 i_329 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [13]), .B1(
      \r_values[1] [6]), .B2(\r_weights[1] [12]), .ZN(n_518));
   AOI21_X1 i_330 (.A(n_519), .B1(n_521), .B2(n_1694), .ZN(n_1693));
   INV_X1 i_331 (.A(n_520), .ZN(n_519));
   OAI21_X1 i_332 (.A(n_1776), .B1(n_522), .B2(n_1694), .ZN(n_520));
   AOI21_X1 i_333 (.A(n_522), .B1(n_1776), .B2(n_521), .ZN(n_1694));
   NAND3_X1 i_334 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [15]), .A3(n_588), 
      .ZN(n_521));
   AOI21_X1 i_335 (.A(n_588), .B1(\r_values[1] [3]), .B2(\r_weights[1] [15]), 
      .ZN(n_522));
   INV_X1 i_336 (.A(n_523), .ZN(n_1595));
   AOI22_X1 i_337 (.A1(\sums[0] [17]), .A2(n_680), .B1(n_591), .B2(n_590), 
      .ZN(n_523));
   OAI21_X1 i_338 (.A(n_526), .B1(n_529), .B2(n_528), .ZN(n_1532));
   OAI21_X1 i_339 (.A(n_533), .B1(n_536), .B2(n_535), .ZN(n_1539));
   OAI21_X1 i_340 (.A(n_542), .B1(n_547), .B2(n_546), .ZN(n_1546));
   OAI21_X1 i_341 (.A(n_549), .B1(n_554), .B2(n_553), .ZN(n_1553));
   AOI21_X1 i_342 (.A(n_560), .B1(n_561), .B2(n_556), .ZN(n_1560));
   OAI22_X1 i_343 (.A1(n_744), .A2(n_566), .B1(n_645), .B2(n_567), .ZN(n_1567));
   OAI22_X1 i_344 (.A1(n_748), .A2(n_576), .B1(n_649), .B2(n_577), .ZN(n_1574));
   OAI22_X1 i_345 (.A1(n_754), .A2(n_582), .B1(n_667), .B2(n_583), .ZN(n_1581));
   OAI21_X1 i_346 (.A(n_587), .B1(n_673), .B2(n_589), .ZN(n_1588));
   XOR2_X1 i_347 (.A(n_529), .B(n_525), .Z(n_1531));
   NAND2_X1 i_348 (.A1(n_527), .A2(n_526), .ZN(n_525));
   NAND3_X1 i_349 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [4]), .A3(n_596), 
      .ZN(n_526));
   INV_X1 i_350 (.A(n_528), .ZN(n_527));
   AOI21_X1 i_351 (.A(n_596), .B1(\r_values[0] [13]), .B2(\r_weights[0] [4]), 
      .ZN(n_528));
   NAND2_X1 i_352 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [2]), .ZN(n_529));
   XOR2_X1 i_353 (.A(n_536), .B(n_532), .Z(n_1538));
   NAND2_X1 i_354 (.A1(n_534), .A2(n_533), .ZN(n_532));
   NAND3_X1 i_355 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [7]), .A3(n_603), 
      .ZN(n_533));
   INV_X1 i_356 (.A(n_535), .ZN(n_534));
   AOI21_X1 i_357 (.A(n_603), .B1(\r_values[0] [10]), .B2(\r_weights[0] [7]), 
      .ZN(n_535));
   NAND2_X1 i_358 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [5]), .ZN(n_536));
   XOR2_X1 i_359 (.A(n_547), .B(n_541), .Z(n_1545));
   NAND2_X1 i_360 (.A1(n_545), .A2(n_542), .ZN(n_541));
   NAND3_X1 i_361 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [10]), .A3(n_621), 
      .ZN(n_542));
   INV_X1 i_362 (.A(n_546), .ZN(n_545));
   AOI21_X1 i_363 (.A(n_621), .B1(\r_values[0] [7]), .B2(\r_weights[0] [10]), 
      .ZN(n_546));
   NAND2_X1 i_364 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [8]), .ZN(n_547));
   XOR2_X1 i_365 (.A(n_554), .B(n_548), .Z(n_1552));
   NAND2_X1 i_366 (.A1(n_552), .A2(n_549), .ZN(n_548));
   NAND3_X1 i_367 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [13]), .A3(n_629), 
      .ZN(n_549));
   INV_X1 i_368 (.A(n_553), .ZN(n_552));
   AOI21_X1 i_369 (.A(n_629), .B1(\r_values[0] [4]), .B2(\r_weights[0] [13]), 
      .ZN(n_553));
   NAND2_X1 i_370 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [11]), .ZN(n_554));
   XOR2_X1 i_371 (.A(n_561), .B(n_555), .Z(n_1559));
   NAND2_X1 i_372 (.A1(n_559), .A2(n_556), .ZN(n_555));
   NAND3_X1 i_373 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [2]), .A3(n_636), 
      .ZN(n_556));
   INV_X1 i_374 (.A(n_560), .ZN(n_559));
   AOI21_X1 i_375 (.A(n_636), .B1(\r_values[1] [15]), .B2(\r_weights[1] [2]), 
      .ZN(n_560));
   NAND2_X1 i_376 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [14]), .ZN(n_561));
   XOR2_X1 i_377 (.A(n_642), .B(n_562), .Z(n_1566));
   AOI21_X1 i_378 (.A(n_567), .B1(n_741), .B2(n_563), .ZN(n_562));
   INV_X1 i_379 (.A(n_566), .ZN(n_563));
   NAND2_X1 i_380 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [5]), .ZN(n_566));
   AOI22_X1 i_381 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [5]), .B1(
      \r_values[1] [13]), .B2(\r_weights[1] [4]), .ZN(n_567));
   XOR2_X1 i_382 (.A(n_648), .B(n_568), .Z(n_1573));
   AOI21_X1 i_383 (.A(n_577), .B1(n_747), .B2(n_569), .ZN(n_568));
   INV_X1 i_384 (.A(n_576), .ZN(n_569));
   NAND2_X1 i_385 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [8]), .ZN(n_576));
   AOI22_X1 i_386 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [8]), .B1(
      \r_values[1] [10]), .B2(\r_weights[1] [7]), .ZN(n_577));
   XOR2_X1 i_387 (.A(n_666), .B(n_580), .Z(n_1580));
   AOI21_X1 i_388 (.A(n_583), .B1(n_753), .B2(n_581), .ZN(n_580));
   INV_X1 i_389 (.A(n_582), .ZN(n_581));
   NAND2_X1 i_390 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [11]), .ZN(n_582));
   AOI22_X1 i_391 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [11]), .B1(
      \r_values[1] [7]), .B2(\r_weights[1] [10]), .ZN(n_583));
   XOR2_X1 i_392 (.A(n_670), .B(n_584), .Z(n_1587));
   AOI21_X1 i_393 (.A(n_589), .B1(n_758), .B2(n_588), .ZN(n_584));
   NAND2_X1 i_394 (.A1(n_758), .A2(n_588), .ZN(n_587));
   AND2_X1 i_395 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [14]), .ZN(n_588));
   AOI22_X1 i_396 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [14]), .B1(
      \r_values[1] [4]), .B2(\r_weights[1] [13]), .ZN(n_589));
   XOR2_X1 i_397 (.A(n_591), .B(n_590), .Z(n_1594));
   OAI21_X1 i_398 (.A(n_677), .B1(n_759), .B2(n_676), .ZN(n_590));
   XNOR2_X1 i_399 (.A(\sums[0] [17]), .B(n_681), .ZN(n_591));
   OAI21_X1 i_400 (.A(n_595), .B1(n_600), .B2(n_598), .ZN(n_1424));
   OAI21_X1 i_401 (.A(n_602), .B1(n_618), .B2(n_615), .ZN(n_1431));
   OAI21_X1 i_402 (.A(n_620), .B1(n_626), .B2(n_625), .ZN(n_1438));
   OAI21_X1 i_403 (.A(n_628), .B1(n_633), .B2(n_632), .ZN(n_1445));
   OAI21_X1 i_404 (.A(n_635), .B1(n_640), .B2(n_639), .ZN(n_1452));
   OAI22_X1 i_405 (.A1(n_827), .A2(n_645), .B1(n_738), .B2(n_646), .ZN(n_1459));
   OAI22_X1 i_406 (.A1(n_855), .A2(n_649), .B1(n_744), .B2(n_662), .ZN(n_1466));
   OAI22_X1 i_407 (.A1(n_861), .A2(n_667), .B1(n_748), .B2(n_668), .ZN(n_1473));
   OAI22_X1 i_408 (.A1(n_867), .A2(n_673), .B1(n_754), .B2(n_674), .ZN(n_1480));
   XOR2_X1 i_409 (.A(n_600), .B(n_594), .Z(n_1423));
   NAND2_X1 i_410 (.A1(n_597), .A2(n_595), .ZN(n_594));
   NAND2_X1 i_411 (.A1(n_787), .A2(n_596), .ZN(n_595));
   AND2_X1 i_412 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [3]), .ZN(n_596));
   INV_X1 i_413 (.A(n_598), .ZN(n_597));
   AOI22_X1 i_414 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [3]), .ZN(n_598));
   NAND2_X1 i_415 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [1]), .ZN(n_600));
   XOR2_X1 i_416 (.A(n_618), .B(n_601), .Z(n_1430));
   NAND2_X1 i_417 (.A1(n_614), .A2(n_602), .ZN(n_601));
   NAND2_X1 i_418 (.A1(n_797), .A2(n_603), .ZN(n_602));
   AND2_X1 i_419 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [6]), .ZN(n_603));
   INV_X1 i_420 (.A(n_615), .ZN(n_614));
   AOI22_X1 i_421 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [6]), .ZN(n_615));
   NAND2_X1 i_422 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [4]), .ZN(n_618));
   XOR2_X1 i_423 (.A(n_626), .B(n_619), .Z(n_1437));
   NAND2_X1 i_424 (.A1(n_622), .A2(n_620), .ZN(n_619));
   NAND2_X1 i_425 (.A1(n_805), .A2(n_621), .ZN(n_620));
   AND2_X1 i_426 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [9]), .ZN(n_621));
   INV_X1 i_427 (.A(n_625), .ZN(n_622));
   AOI22_X1 i_428 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [9]), .ZN(n_625));
   NAND2_X1 i_429 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [7]), .ZN(n_626));
   XOR2_X1 i_430 (.A(n_633), .B(n_627), .Z(n_1444));
   NAND2_X1 i_431 (.A1(n_631), .A2(n_628), .ZN(n_627));
   NAND2_X1 i_432 (.A1(n_812), .A2(n_629), .ZN(n_628));
   AND2_X1 i_433 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [12]), .ZN(n_629));
   INV_X1 i_434 (.A(n_632), .ZN(n_631));
   AOI22_X1 i_435 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [11]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [12]), .ZN(n_632));
   NAND2_X1 i_436 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [10]), .ZN(n_633));
   XOR2_X1 i_437 (.A(n_640), .B(n_634), .Z(n_1451));
   NAND2_X1 i_438 (.A1(n_638), .A2(n_635), .ZN(n_634));
   NAND2_X1 i_439 (.A1(n_819), .A2(n_636), .ZN(n_635));
   AND2_X1 i_440 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [15]), .ZN(n_636));
   INV_X1 i_441 (.A(n_639), .ZN(n_638));
   AOI22_X1 i_442 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [14]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [15]), .ZN(n_639));
   NAND2_X1 i_443 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [13]), .ZN(n_640));
   XOR2_X1 i_444 (.A(n_737), .B(n_641), .Z(n_1458));
   AOI21_X1 i_445 (.A(n_646), .B1(n_826), .B2(n_642), .ZN(n_641));
   INV_X1 i_446 (.A(n_645), .ZN(n_642));
   NAND2_X1 i_447 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [3]), .ZN(n_645));
   AOI22_X1 i_448 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [3]), .B1(
      \r_values[1] [14]), .B2(\r_weights[1] [2]), .ZN(n_646));
   XOR2_X1 i_449 (.A(n_741), .B(n_647), .Z(n_1465));
   AOI21_X1 i_450 (.A(n_662), .B1(n_854), .B2(n_648), .ZN(n_647));
   INV_X1 i_451 (.A(n_649), .ZN(n_648));
   NAND2_X1 i_452 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [6]), .ZN(n_649));
   AOI22_X1 i_453 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [6]), .B1(
      \r_values[1] [11]), .B2(\r_weights[1] [5]), .ZN(n_662));
   XOR2_X1 i_454 (.A(n_747), .B(n_663), .Z(n_1472));
   AOI21_X1 i_455 (.A(n_668), .B1(n_860), .B2(n_666), .ZN(n_663));
   INV_X1 i_456 (.A(n_667), .ZN(n_666));
   NAND2_X1 i_457 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [9]), .ZN(n_667));
   AOI22_X1 i_458 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [9]), .B1(
      \r_values[1] [8]), .B2(\r_weights[1] [8]), .ZN(n_668));
   XOR2_X1 i_459 (.A(n_753), .B(n_669), .Z(n_1479));
   AOI21_X1 i_460 (.A(n_674), .B1(n_864), .B2(n_670), .ZN(n_669));
   INV_X1 i_461 (.A(n_673), .ZN(n_670));
   NAND2_X1 i_462 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [12]), .ZN(n_673));
   AOI22_X1 i_463 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [12]), .B1(
      \r_values[1] [5]), .B2(\r_weights[1] [11]), .ZN(n_674));
   XOR2_X1 i_464 (.A(n_758), .B(n_675), .Z(n_1486));
   AOI21_X1 i_465 (.A(n_676), .B1(n_871), .B2(n_680), .ZN(n_675));
   AOI22_X1 i_466 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [15]), .B1(
      \r_values[1] [2]), .B2(\r_weights[1] [14]), .ZN(n_676));
   NAND2_X1 i_467 (.A1(n_871), .A2(n_680), .ZN(n_677));
   INV_X1 i_468 (.A(n_681), .ZN(n_680));
   NAND2_X1 i_469 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [15]), .ZN(n_681));
   OAI21_X1 i_470 (.A(n_683), .B1(n_688), .B2(n_687), .ZN(n_1310));
   OAI21_X1 i_471 (.A(n_690), .B1(n_695), .B2(n_694), .ZN(n_1317));
   OAI21_X1 i_472 (.A(n_697), .B1(n_702), .B2(n_701), .ZN(n_1324));
   OAI21_X1 i_473 (.A(n_704), .B1(n_723), .B2(n_720), .ZN(n_1331));
   OAI21_X1 i_474 (.A(n_725), .B1(n_730), .B2(n_727), .ZN(n_1338));
   AOI21_X1 i_475 (.A(n_733), .B1(n_739), .B2(n_734), .ZN(n_1345));
   OAI22_X1 i_476 (.A1(n_942), .A2(n_744), .B1(n_827), .B2(n_745), .ZN(n_1352));
   OAI22_X1 i_477 (.A1(n_948), .A2(n_748), .B1(n_855), .B2(n_751), .ZN(n_1359));
   OAI22_X1 i_478 (.A1(n_954), .A2(n_754), .B1(n_861), .B2(n_755), .ZN(n_1366));
   OAI22_X1 i_479 (.A1(n_961), .A2(n_759), .B1(n_867), .B2(n_760), .ZN(n_1373));
   XOR2_X1 i_480 (.A(n_688), .B(n_682), .Z(n_1309));
   NAND2_X1 i_481 (.A1(n_684), .A2(n_683), .ZN(n_682));
   NAND3_X1 i_482 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [1]), .A3(n_787), 
      .ZN(n_683));
   INV_X1 i_483 (.A(n_687), .ZN(n_684));
   AOI21_X1 i_484 (.A(n_787), .B1(\r_values[0] [14]), .B2(\r_weights[0] [1]), 
      .ZN(n_687));
   NAND2_X1 i_485 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [0]), .ZN(n_688));
   XOR2_X1 i_486 (.A(n_695), .B(n_689), .Z(n_1316));
   NAND2_X1 i_487 (.A1(n_691), .A2(n_690), .ZN(n_689));
   NAND3_X1 i_488 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [4]), .A3(n_797), 
      .ZN(n_690));
   INV_X1 i_489 (.A(n_694), .ZN(n_691));
   AOI21_X1 i_490 (.A(n_797), .B1(\r_values[0] [11]), .B2(\r_weights[0] [4]), 
      .ZN(n_694));
   NAND2_X1 i_491 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [3]), .ZN(n_695));
   XOR2_X1 i_492 (.A(n_702), .B(n_696), .Z(n_1323));
   NAND2_X1 i_493 (.A1(n_698), .A2(n_697), .ZN(n_696));
   NAND3_X1 i_494 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [7]), .A3(n_805), 
      .ZN(n_697));
   INV_X1 i_495 (.A(n_701), .ZN(n_698));
   AOI21_X1 i_496 (.A(n_805), .B1(\r_values[0] [8]), .B2(\r_weights[0] [7]), 
      .ZN(n_701));
   NAND2_X1 i_497 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [6]), .ZN(n_702));
   XOR2_X1 i_498 (.A(n_723), .B(n_703), .Z(n_1330));
   NAND2_X1 i_499 (.A1(n_719), .A2(n_704), .ZN(n_703));
   NAND3_X1 i_500 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [10]), .A3(n_812), 
      .ZN(n_704));
   INV_X1 i_501 (.A(n_720), .ZN(n_719));
   AOI21_X1 i_502 (.A(n_812), .B1(\r_values[0] [5]), .B2(\r_weights[0] [10]), 
      .ZN(n_720));
   NAND2_X1 i_503 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [9]), .ZN(n_723));
   XOR2_X1 i_504 (.A(n_730), .B(n_724), .Z(n_1337));
   NAND2_X1 i_505 (.A1(n_726), .A2(n_725), .ZN(n_724));
   NAND3_X1 i_506 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [13]), .A3(n_819), 
      .ZN(n_725));
   INV_X1 i_507 (.A(n_727), .ZN(n_726));
   AOI21_X1 i_508 (.A(n_819), .B1(\r_values[0] [2]), .B2(\r_weights[0] [13]), 
      .ZN(n_727));
   NAND2_X1 i_509 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [12]), .ZN(n_730));
   XOR2_X1 i_510 (.A(n_739), .B(n_731), .Z(n_1344));
   NAND2_X1 i_511 (.A1(n_734), .A2(n_732), .ZN(n_731));
   INV_X1 i_512 (.A(n_733), .ZN(n_732));
   AOI22_X1 i_514 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [1]), .B1(
      \r_values[1] [15]), .B2(\r_weights[1] [0]), .ZN(n_733));
   NAND2_X1 i_515 (.A1(n_849), .A2(n_737), .ZN(n_734));
   INV_X1 i_516 (.A(n_738), .ZN(n_737));
   NAND2_X1 i_517 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [1]), .ZN(n_738));
   NAND2_X1 i_518 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [15]), .ZN(n_739));
   XOR2_X1 i_519 (.A(n_826), .B(n_740), .Z(n_1351));
   AOI21_X1 i_520 (.A(n_745), .B1(n_941), .B2(n_741), .ZN(n_740));
   INV_X1 i_521 (.A(n_744), .ZN(n_741));
   NAND2_X1 i_522 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [4]), .ZN(n_744));
   AOI22_X1 i_523 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [4]), .B1(
      \r_values[1] [12]), .B2(\r_weights[1] [3]), .ZN(n_745));
   XOR2_X1 i_524 (.A(n_854), .B(n_746), .Z(n_1358));
   AOI21_X1 i_525 (.A(n_751), .B1(n_947), .B2(n_747), .ZN(n_746));
   INV_X1 i_526 (.A(n_748), .ZN(n_747));
   NAND2_X1 i_527 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [7]), .ZN(n_748));
   AOI22_X1 i_528 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [7]), .B1(
      \r_values[1] [9]), .B2(\r_weights[1] [6]), .ZN(n_751));
   XOR2_X1 i_529 (.A(n_860), .B(n_752), .Z(n_1365));
   AOI21_X1 i_530 (.A(n_755), .B1(n_953), .B2(n_753), .ZN(n_752));
   INV_X1 i_531 (.A(n_754), .ZN(n_753));
   NAND2_X1 i_532 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [10]), .ZN(n_754));
   AOI22_X1 i_533 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [10]), .B1(
      \r_values[1] [6]), .B2(\r_weights[1] [9]), .ZN(n_755));
   XOR2_X1 i_534 (.A(n_864), .B(n_757), .Z(n_1372));
   AOI21_X1 i_535 (.A(n_760), .B1(n_960), .B2(n_758), .ZN(n_757));
   INV_X1 i_538 (.A(n_759), .ZN(n_758));
   NAND2_X1 i_539 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [13]), .ZN(n_759));
   AOI22_X1 i_540 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [13]), .B1(
      \r_values[1] [3]), .B2(\r_weights[1] [12]), .ZN(n_760));
   AOI21_X1 i_541 (.A(n_779), .B1(n_783), .B2(n_1379), .ZN(n_1378));
   INV_X1 i_542 (.A(n_780), .ZN(n_779));
   OAI21_X1 i_543 (.A(n_1775), .B1(n_784), .B2(n_1379), .ZN(n_780));
   AOI21_X1 i_544 (.A(n_784), .B1(n_1775), .B2(n_783), .ZN(n_1379));
   NAND3_X1 i_545 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [15]), .A3(n_871), 
      .ZN(n_783));
   AOI21_X1 i_546 (.A(n_871), .B1(\r_values[1] [0]), .B2(\r_weights[1] [15]), 
      .ZN(n_784));
   OAI21_X1 i_547 (.A(n_786), .B1(n_792), .B2(n_791), .ZN(n_1206));
   OAI21_X1 i_548 (.A(n_794), .B1(n_800), .B2(n_799), .ZN(n_1213));
   OAI21_X1 i_549 (.A(n_804), .B1(n_808), .B2(n_807), .ZN(n_1220));
   OAI21_X1 i_550 (.A(n_811), .B1(n_815), .B2(n_814), .ZN(n_1227));
   OAI21_X1 i_551 (.A(n_818), .B1(n_824), .B2(n_821), .ZN(n_1234));
   OAI22_X1 i_552 (.A1(n_1029), .A2(n_827), .B1(n_850), .B2(n_828), .ZN(n_1241));
   OAI22_X1 i_553 (.A1(n_1035), .A2(n_855), .B1(n_942), .B2(n_856), .ZN(n_1248));
   OAI22_X1 i_554 (.A1(n_1039), .A2(n_861), .B1(n_948), .B2(n_862), .ZN(n_1255));
   OAI22_X1 i_555 (.A1(n_1045), .A2(n_867), .B1(n_954), .B2(n_868), .ZN(n_1262));
   OAI21_X1 i_556 (.A(n_870), .B1(n_961), .B2(n_874), .ZN(n_1269));
   XOR2_X1 i_557 (.A(n_792), .B(n_785), .Z(n_1205));
   NAND2_X1 i_558 (.A1(n_790), .A2(n_786), .ZN(n_785));
   NAND2_X1 i_559 (.A1(n_882), .A2(n_787), .ZN(n_786));
   AND2_X1 i_560 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [2]), .ZN(n_787));
   INV_X1 i_561 (.A(n_791), .ZN(n_790));
   AOI22_X1 i_562 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [13]), .B2(\r_weights[0] [1]), .ZN(n_791));
   NAND2_X1 i_563 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [0]), .ZN(n_792));
   XOR2_X1 i_564 (.A(n_800), .B(n_793), .Z(n_1212));
   NAND2_X1 i_565 (.A1(n_798), .A2(n_794), .ZN(n_793));
   NAND2_X1 i_566 (.A1(n_890), .A2(n_797), .ZN(n_794));
   AND2_X1 i_570 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [5]), .ZN(n_797));
   INV_X1 i_571 (.A(n_799), .ZN(n_798));
   AOI22_X1 i_572 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [4]), .ZN(n_799));
   NAND2_X1 i_573 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [3]), .ZN(n_800));
   XOR2_X1 i_574 (.A(n_808), .B(n_801), .Z(n_1219));
   NAND2_X1 i_575 (.A1(n_806), .A2(n_804), .ZN(n_801));
   NAND2_X1 i_576 (.A1(n_898), .A2(n_805), .ZN(n_804));
   AND2_X1 i_577 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [8]), .ZN(n_805));
   INV_X1 i_578 (.A(n_807), .ZN(n_806));
   AOI22_X1 i_579 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [7]), .ZN(n_807));
   NAND2_X1 i_580 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [6]), .ZN(n_808));
   XOR2_X1 i_581 (.A(n_815), .B(n_810), .Z(n_1226));
   NAND2_X1 i_582 (.A1(n_813), .A2(n_811), .ZN(n_810));
   NAND2_X1 i_583 (.A1(n_928), .A2(n_812), .ZN(n_811));
   AND2_X1 i_584 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [11]), .ZN(n_812));
   INV_X1 i_585 (.A(n_814), .ZN(n_813));
   AOI22_X1 i_586 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [11]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [10]), .ZN(n_814));
   NAND2_X1 i_587 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [9]), .ZN(n_815));
   XOR2_X1 i_588 (.A(n_824), .B(n_817), .Z(n_1233));
   NAND2_X1 i_589 (.A1(n_820), .A2(n_818), .ZN(n_817));
   NAND2_X1 i_590 (.A1(n_936), .A2(n_819), .ZN(n_818));
   AND2_X1 i_591 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [14]), .ZN(n_819));
   INV_X1 i_592 (.A(n_821), .ZN(n_820));
   AOI22_X1 i_593 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [14]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [13]), .ZN(n_821));
   NAND2_X1 i_594 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [12]), .ZN(n_824));
   XOR2_X1 i_595 (.A(n_849), .B(n_825), .Z(n_1240));
   AOI21_X1 i_596 (.A(n_828), .B1(n_1028), .B2(n_826), .ZN(n_825));
   INV_X1 i_597 (.A(n_827), .ZN(n_826));
   NAND2_X1 i_603 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [2]), .ZN(n_827));
   AOI22_X1 i_604 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [2]), .B1(
      \r_values[1] [13]), .B2(\r_weights[1] [1]), .ZN(n_828));
   INV_X1 i_605 (.A(n_850), .ZN(n_849));
   NAND2_X1 i_606 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [0]), .ZN(n_850));
   XOR2_X1 i_607 (.A(n_941), .B(n_853), .Z(n_1247));
   AOI21_X1 i_608 (.A(n_856), .B1(n_1032), .B2(n_854), .ZN(n_853));
   INV_X1 i_609 (.A(n_855), .ZN(n_854));
   NAND2_X1 i_610 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [5]), .ZN(n_855));
   AOI22_X1 i_611 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [5]), .B1(
      \r_values[1] [10]), .B2(\r_weights[1] [4]), .ZN(n_856));
   XOR2_X1 i_612 (.A(n_947), .B(n_857), .Z(n_1254));
   AOI21_X1 i_613 (.A(n_862), .B1(n_1038), .B2(n_860), .ZN(n_857));
   INV_X1 i_614 (.A(n_861), .ZN(n_860));
   NAND2_X1 i_615 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [8]), .ZN(n_861));
   AOI22_X1 i_616 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [8]), .B1(
      \r_values[1] [7]), .B2(\r_weights[1] [7]), .ZN(n_862));
   XOR2_X1 i_617 (.A(n_953), .B(n_863), .Z(n_1261));
   AOI21_X1 i_618 (.A(n_868), .B1(n_1044), .B2(n_864), .ZN(n_863));
   INV_X1 i_619 (.A(n_867), .ZN(n_864));
   NAND2_X1 i_620 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [11]), .ZN(n_867));
   AOI22_X1 i_621 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [11]), .B1(
      \r_values[1] [4]), .B2(\r_weights[1] [10]), .ZN(n_868));
   XOR2_X1 i_622 (.A(n_960), .B(n_869), .Z(n_1268));
   AOI21_X1 i_623 (.A(n_874), .B1(n_964), .B2(n_871), .ZN(n_869));
   NAND2_X1 i_624 (.A1(n_964), .A2(n_871), .ZN(n_870));
   AND2_X1 i_625 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [14]), .ZN(n_871));
   AOI22_X1 i_626 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [14]), .B1(
      \r_values[1] [1]), .B2(\r_weights[1] [13]), .ZN(n_874));
   OAI21_X1 i_627 (.A(n_875), .B1(n_1772), .B2(n_967), .ZN(n_1168));
   OAI21_X1 i_628 (.A(n_1051), .B1(\sums[0] [13]), .B2(n_964), .ZN(n_875));
   OAI21_X1 i_629 (.A(n_877), .B1(n_883), .B2(n_881), .ZN(n_1105));
   OAI21_X1 i_630 (.A(n_885), .B1(n_891), .B2(n_889), .ZN(n_1112));
   OAI21_X1 i_631 (.A(n_895), .B1(n_899), .B2(n_897), .ZN(n_1119));
   OAI21_X1 i_632 (.A(n_903), .B1(n_929), .B2(n_905), .ZN(n_1126));
   AOI21_X1 i_633 (.A(n_935), .B1(n_939), .B2(n_933), .ZN(n_1133));
   OAI22_X1 i_634 (.A1(n_1114), .A2(n_942), .B1(n_1029), .B2(n_943), .ZN(n_1140));
   OAI22_X1 i_635 (.A1(n_1122), .A2(n_948), .B1(n_1035), .B2(n_949), .ZN(n_1147));
   OAI22_X1 i_636 (.A1(n_1128), .A2(n_954), .B1(n_1039), .B2(n_955), .ZN(n_1154));
   OAI21_X1 i_637 (.A(n_957), .B1(n_1045), .B2(n_962), .ZN(n_1161));
   XOR2_X1 i_638 (.A(n_883), .B(n_876), .Z(n_1104));
   NAND2_X1 i_645 (.A1(n_878), .A2(n_877), .ZN(n_876));
   NAND3_X1 i_646 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [2]), .A3(n_882), 
      .ZN(n_877));
   INV_X1 i_647 (.A(n_881), .ZN(n_878));
   AOI21_X1 i_648 (.A(n_882), .B1(\r_values[0] [11]), .B2(\r_weights[0] [2]), 
      .ZN(n_881));
   AND2_X1 i_649 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [1]), .ZN(n_882));
   NAND2_X1 i_650 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [0]), .ZN(n_883));
   XOR2_X1 i_651 (.A(n_891), .B(n_884), .Z(n_1111));
   NAND2_X1 i_652 (.A1(n_888), .A2(n_885), .ZN(n_884));
   NAND3_X1 i_653 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [5]), .A3(n_890), 
      .ZN(n_885));
   INV_X1 i_654 (.A(n_889), .ZN(n_888));
   AOI21_X1 i_655 (.A(n_890), .B1(\r_values[0] [8]), .B2(\r_weights[0] [5]), 
      .ZN(n_889));
   AND2_X1 i_656 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [4]), .ZN(n_890));
   NAND2_X1 i_657 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [3]), .ZN(n_891));
   XOR2_X1 i_658 (.A(n_899), .B(n_892), .Z(n_1118));
   NAND2_X1 i_659 (.A1(n_896), .A2(n_895), .ZN(n_892));
   NAND3_X1 i_660 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [8]), .A3(n_898), 
      .ZN(n_895));
   INV_X1 i_661 (.A(n_897), .ZN(n_896));
   AOI21_X1 i_662 (.A(n_898), .B1(\r_values[0] [5]), .B2(\r_weights[0] [8]), 
      .ZN(n_897));
   AND2_X1 i_663 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [7]), .ZN(n_898));
   NAND2_X1 i_664 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [6]), .ZN(n_899));
   XOR2_X1 i_665 (.A(n_929), .B(n_902), .Z(n_1125));
   NAND2_X1 i_666 (.A1(n_904), .A2(n_903), .ZN(n_902));
   NAND3_X1 i_667 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [11]), .A3(n_928), 
      .ZN(n_903));
   INV_X1 i_668 (.A(n_905), .ZN(n_904));
   AOI21_X1 i_669 (.A(n_928), .B1(\r_values[0] [2]), .B2(\r_weights[0] [11]), 
      .ZN(n_905));
   AND2_X1 i_670 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [10]), .ZN(n_928));
   NAND2_X1 i_671 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [9]), .ZN(n_929));
   XOR2_X1 i_672 (.A(n_939), .B(n_932), .Z(n_1132));
   NAND2_X1 i_673 (.A1(n_934), .A2(n_933), .ZN(n_932));
   NAND3_X1 i_674 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [0]), .A3(n_936), 
      .ZN(n_933));
   INV_X1 i_675 (.A(n_935), .ZN(n_934));
   AOI21_X1 i_676 (.A(n_936), .B1(\r_values[1] [13]), .B2(\r_weights[1] [0]), 
      .ZN(n_935));
   AND2_X1 i_677 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [13]), .ZN(n_936));
   NAND2_X1 i_678 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [12]), .ZN(n_939));
   XOR2_X1 i_679 (.A(n_1028), .B(n_940), .Z(n_1139));
   AOI21_X1 i_680 (.A(n_943), .B1(n_1113), .B2(n_941), .ZN(n_940));
   INV_X1 i_681 (.A(n_942), .ZN(n_941));
   NAND2_X1 i_682 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [3]), .ZN(n_942));
   AOI22_X1 i_683 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [3]), .B1(
      \r_values[1] [11]), .B2(\r_weights[1] [2]), .ZN(n_943));
   XOR2_X1 i_684 (.A(n_1032), .B(n_946), .Z(n_1146));
   AOI21_X1 i_685 (.A(n_949), .B1(n_1121), .B2(n_947), .ZN(n_946));
   INV_X1 i_686 (.A(n_948), .ZN(n_947));
   NAND2_X1 i_687 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [6]), .ZN(n_948));
   AOI22_X1 i_695 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [6]), .B1(
      \r_values[1] [8]), .B2(\r_weights[1] [5]), .ZN(n_949));
   XOR2_X1 i_696 (.A(n_1038), .B(n_950), .Z(n_1153));
   AOI21_X1 i_697 (.A(n_955), .B1(n_1127), .B2(n_953), .ZN(n_950));
   INV_X1 i_698 (.A(n_954), .ZN(n_953));
   NAND2_X1 i_699 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [9]), .ZN(n_954));
   AOI22_X1 i_700 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [9]), .B1(
      \r_values[1] [5]), .B2(\r_weights[1] [8]), .ZN(n_955));
   XOR2_X1 i_701 (.A(n_1044), .B(n_956), .Z(n_1160));
   AOI21_X1 i_702 (.A(n_962), .B1(n_1134), .B2(n_960), .ZN(n_956));
   NAND2_X1 i_703 (.A1(n_1134), .A2(n_960), .ZN(n_957));
   INV_X1 i_704 (.A(n_961), .ZN(n_960));
   NAND2_X1 i_705 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [12]), .ZN(n_961));
   AOI22_X1 i_706 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [12]), .B1(
      \r_values[1] [2]), .B2(\r_weights[1] [11]), .ZN(n_962));
   XNOR2_X1 i_707 (.A(n_1051), .B(n_963), .ZN(n_1167));
   OAI22_X1 i_708 (.A1(n_1772), .A2(n_967), .B1(\sums[0] [13]), .B2(n_964), 
      .ZN(n_963));
   INV_X1 i_709 (.A(n_967), .ZN(n_964));
   NAND2_X1 i_710 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [13]), .ZN(n_967));
   OAI21_X1 i_711 (.A(n_969), .B1(n_974), .B2(n_971), .ZN(n_1013));
   OAI21_X1 i_712 (.A(n_976), .B1(n_981), .B2(n_978), .ZN(n_1020));
   OAI21_X1 i_713 (.A(n_983), .B1(n_1014), .B2(n_1011), .ZN(n_1027));
   OAI21_X1 i_714 (.A(n_1016), .B1(n_1021), .B2(n_1018), .ZN(n_1034));
   AOI21_X1 i_715 (.A(n_1024), .B1(n_1030), .B2(n_1025), .ZN(n_1041));
   OAI22_X1 i_716 (.A1(n_1209), .A2(n_1035), .B1(n_1114), .B2(n_1036), .ZN(
      n_1048));
   OAI22_X1 i_717 (.A1(n_1216), .A2(n_1039), .B1(n_1122), .B2(n_1042), .ZN(
      n_1055));
   OAI22_X1 i_718 (.A1(n_1222), .A2(n_1045), .B1(n_1128), .B2(n_1046), .ZN(
      n_1062));
   XOR2_X1 i_719 (.A(n_974), .B(n_968), .Z(n_1012));
   NAND2_X1 i_720 (.A1(n_970), .A2(n_969), .ZN(n_968));
   NAND4_X1 i_721 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [11]), .A4(\r_weights[0] [1]), .ZN(n_969));
   INV_X1 i_722 (.A(n_971), .ZN(n_970));
   AOI22_X1 i_723 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [11]), .B2(\r_weights[0] [1]), .ZN(n_971));
   NAND2_X1 i_724 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [0]), .ZN(n_974));
   XOR2_X1 i_725 (.A(n_981), .B(n_975), .Z(n_1019));
   NAND2_X1 i_726 (.A1(n_977), .A2(n_976), .ZN(n_975));
   NAND4_X1 i_727 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [8]), .A4(\r_weights[0] [4]), .ZN(n_976));
   INV_X1 i_728 (.A(n_978), .ZN(n_977));
   AOI22_X1 i_729 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [8]), .B2(\r_weights[0] [4]), .ZN(n_978));
   NAND2_X1 i_730 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [3]), .ZN(n_981));
   XOR2_X1 i_731 (.A(n_1014), .B(n_982), .Z(n_1026));
   NAND2_X1 i_732 (.A1(n_1010), .A2(n_983), .ZN(n_982));
   NAND4_X1 i_733 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [8]), .A3(
      \r_values[0] [5]), .A4(\r_weights[0] [7]), .ZN(n_983));
   INV_X1 i_734 (.A(n_1011), .ZN(n_1010));
   AOI22_X1 i_735 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [5]), .B2(\r_weights[0] [7]), .ZN(n_1011));
   NAND2_X1 i_736 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [6]), .ZN(n_1014));
   XOR2_X1 i_746 (.A(n_1021), .B(n_1015), .Z(n_1033));
   NAND2_X1 i_747 (.A1(n_1017), .A2(n_1016), .ZN(n_1015));
   NAND3_X1 i_748 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [10]), .A3(n_1106), 
      .ZN(n_1016));
   INV_X1 i_749 (.A(n_1018), .ZN(n_1017));
   AOI21_X1 i_750 (.A(n_1106), .B1(\r_values[0] [2]), .B2(\r_weights[0] [10]), 
      .ZN(n_1018));
   NAND2_X1 i_751 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [9]), .ZN(n_1021));
   XOR2_X1 i_752 (.A(n_1030), .B(n_1022), .Z(n_1040));
   NAND2_X1 i_753 (.A1(n_1025), .A2(n_1023), .ZN(n_1022));
   INV_X1 i_754 (.A(n_1024), .ZN(n_1023));
   AOI22_X1 i_755 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [1]), .B1(
      \r_values[1] [12]), .B2(\r_weights[1] [0]), .ZN(n_1024));
   NAND2_X1 i_756 (.A1(n_1116), .A2(n_1028), .ZN(n_1025));
   INV_X1 i_757 (.A(n_1029), .ZN(n_1028));
   NAND2_X1 i_758 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [1]), .ZN(n_1029));
   NAND2_X1 i_759 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [12]), .ZN(n_1030));
   XOR2_X1 i_760 (.A(n_1113), .B(n_1031), .Z(n_1047));
   AOI21_X1 i_761 (.A(n_1036), .B1(n_1208), .B2(n_1032), .ZN(n_1031));
   INV_X1 i_762 (.A(n_1035), .ZN(n_1032));
   NAND2_X1 i_763 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [4]), .ZN(n_1035));
   AOI22_X1 i_764 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [4]), .B1(
      \r_values[1] [9]), .B2(\r_weights[1] [3]), .ZN(n_1036));
   XOR2_X1 i_765 (.A(n_1121), .B(n_1037), .Z(n_1054));
   AOI21_X1 i_766 (.A(n_1042), .B1(n_1215), .B2(n_1038), .ZN(n_1037));
   INV_X1 i_767 (.A(n_1039), .ZN(n_1038));
   NAND2_X1 i_768 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [7]), .ZN(n_1039));
   AOI22_X1 i_769 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [7]), .B1(
      \r_values[1] [6]), .B2(\r_weights[1] [6]), .ZN(n_1042));
   XOR2_X1 i_770 (.A(n_1127), .B(n_1043), .Z(n_1061));
   AOI21_X1 i_771 (.A(n_1046), .B1(n_1221), .B2(n_1044), .ZN(n_1043));
   INV_X1 i_772 (.A(n_1045), .ZN(n_1044));
   NAND2_X1 i_773 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [10]), .ZN(n_1045));
   AOI22_X1 i_774 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [10]), .B1(
      \r_values[1] [3]), .B2(\r_weights[1] [9]), .ZN(n_1046));
   AOI21_X1 i_775 (.A(n_1049), .B1(n_1771), .B2(n_1053), .ZN(n_1067));
   INV_X1 i_776 (.A(n_1050), .ZN(n_1049));
   OAI21_X1 i_777 (.A(n_1051), .B1(n_1771), .B2(n_1052), .ZN(n_1050));
   AOI21_X1 i_778 (.A(n_1053), .B1(n_1771), .B2(n_1052), .ZN(n_1051));
   NAND3_X1 i_779 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [12]), .A3(n_1134), 
      .ZN(n_1052));
   AOI21_X1 i_780 (.A(n_1134), .B1(\r_values[1] [0]), .B2(\r_weights[1] [12]), 
      .ZN(n_1053));
   OAI21_X1 i_781 (.A(n_1057), .B1(n_1060), .B2(n_1059), .ZN(n_931));
   OAI21_X1 i_782 (.A(n_1064), .B1(n_1068), .B2(n_1066), .ZN(n_938));
   OAI21_X1 i_783 (.A(n_1070), .B1(n_1073), .B2(n_1072), .ZN(n_945));
   OAI21_X1 i_784 (.A(n_1103), .B1(n_1109), .B2(n_1108), .ZN(n_952));
   OAI22_X1 i_785 (.A1(n_1253), .A2(n_1114), .B1(n_1117), .B2(n_1115), .ZN(n_959));
   OAI22_X1 i_786 (.A1(n_1264), .A2(n_1122), .B1(n_1209), .B2(n_1123), .ZN(n_966));
   OAI22_X1 i_787 (.A1(n_1272), .A2(n_1128), .B1(n_1216), .B2(n_1129), .ZN(n_973));
   OAI21_X1 i_788 (.A(n_1131), .B1(n_1222), .B2(n_1136), .ZN(n_980));
   XOR2_X1 i_789 (.A(n_1060), .B(n_1056), .Z(n_930));
   NAND2_X1 i_790 (.A1(n_1058), .A2(n_1057), .ZN(n_1056));
   NAND4_X1 i_791 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [10]), .A4(\r_weights[0] [1]), .ZN(n_1057));
   INV_X1 i_792 (.A(n_1059), .ZN(n_1058));
   AOI22_X1 i_793 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [10]), .B2(\r_weights[0] [1]), .ZN(n_1059));
   NAND2_X1 i_794 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [0]), .ZN(n_1060));
   XOR2_X1 i_795 (.A(n_1068), .B(n_1063), .Z(n_937));
   NAND2_X1 i_806 (.A1(n_1065), .A2(n_1064), .ZN(n_1063));
   NAND4_X1 i_807 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [7]), .A4(\r_weights[0] [4]), .ZN(n_1064));
   INV_X1 i_808 (.A(n_1066), .ZN(n_1065));
   AOI22_X1 i_809 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [4]), .ZN(n_1066));
   NAND2_X1 i_810 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [3]), .ZN(n_1068));
   XOR2_X1 i_811 (.A(n_1073), .B(n_1069), .Z(n_944));
   NAND2_X1 i_812 (.A1(n_1071), .A2(n_1070), .ZN(n_1069));
   NAND4_X1 i_813 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [8]), .A3(
      \r_values[0] [4]), .A4(\r_weights[0] [7]), .ZN(n_1070));
   INV_X1 i_814 (.A(n_1072), .ZN(n_1071));
   AOI22_X1 i_815 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [7]), .ZN(n_1072));
   NAND2_X1 i_816 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [6]), .ZN(n_1073));
   XOR2_X1 i_817 (.A(n_1109), .B(n_1102), .Z(n_951));
   NAND2_X1 i_818 (.A1(n_1107), .A2(n_1103), .ZN(n_1102));
   NAND2_X1 i_819 (.A1(n_1172), .A2(n_1106), .ZN(n_1103));
   AND2_X1 i_820 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [11]), .ZN(n_1106));
   INV_X1 i_821 (.A(n_1108), .ZN(n_1107));
   AOI22_X1 i_822 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [11]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [10]), .ZN(n_1108));
   NAND2_X1 i_823 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [9]), .ZN(n_1109));
   XOR2_X1 i_824 (.A(n_1116), .B(n_1110), .Z(n_958));
   AOI21_X1 i_825 (.A(n_1115), .B1(n_1252), .B2(n_1113), .ZN(n_1110));
   INV_X1 i_826 (.A(n_1114), .ZN(n_1113));
   NAND2_X1 i_827 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [2]), .ZN(n_1114));
   AOI22_X1 i_828 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [2]), .B1(
      \r_values[1] [10]), .B2(\r_weights[1] [1]), .ZN(n_1115));
   INV_X1 i_829 (.A(n_1117), .ZN(n_1116));
   NAND2_X1 i_830 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [0]), .ZN(n_1117));
   XOR2_X1 i_831 (.A(n_1208), .B(n_1120), .Z(n_965));
   AOI21_X1 i_832 (.A(n_1123), .B1(n_1263), .B2(n_1121), .ZN(n_1120));
   INV_X1 i_833 (.A(n_1122), .ZN(n_1121));
   NAND2_X1 i_834 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [5]), .ZN(n_1122));
   AOI22_X1 i_835 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [5]), .B1(
      \r_values[1] [7]), .B2(\r_weights[1] [4]), .ZN(n_1123));
   XOR2_X1 i_836 (.A(n_1215), .B(n_1124), .Z(n_972));
   AOI21_X1 i_837 (.A(n_1129), .B1(n_1271), .B2(n_1127), .ZN(n_1124));
   INV_X1 i_838 (.A(n_1128), .ZN(n_1127));
   NAND2_X1 i_839 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [8]), .ZN(n_1128));
   AOI22_X1 i_840 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [8]), .B1(
      \r_values[1] [4]), .B2(\r_weights[1] [7]), .ZN(n_1129));
   XNOR2_X1 i_841 (.A(n_1221), .B(n_1130), .ZN(n_979));
   NAND2_X1 i_842 (.A1(n_1135), .A2(n_1131), .ZN(n_1130));
   NAND3_X1 i_843 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [10]), .A3(n_1134), 
      .ZN(n_1131));
   AND2_X1 i_844 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [11]), .ZN(n_1134));
   INV_X1 i_845 (.A(n_1136), .ZN(n_1135));
   AOI22_X1 i_846 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [11]), .B1(
      \r_values[1] [1]), .B2(\r_weights[1] [10]), .ZN(n_1136));
   AOI22_X1 i_847 (.A1(n_1143), .A2(n_1142), .B1(n_1144), .B2(n_1141), .ZN(n_901));
   OAI21_X1 i_848 (.A(n_1148), .B1(n_1151), .B2(n_1150), .ZN(n_852));
   OAI21_X1 i_849 (.A(n_1155), .B1(n_1158), .B2(n_1157), .ZN(n_859));
   OAI21_X1 i_850 (.A(n_1162), .B1(n_1165), .B2(n_1164), .ZN(n_866));
   AOI21_X1 i_851 (.A(n_1171), .B1(n_1203), .B2(n_1169), .ZN(n_873));
   OAI21_X1 i_852 (.A(n_1207), .B1(n_1253), .B2(n_1210), .ZN(n_880));
   OAI21_X1 i_853 (.A(n_1214), .B1(n_1264), .B2(n_1217), .ZN(n_887));
   OAI22_X1 i_854 (.A1(n_1354), .A2(n_1222), .B1(n_1272), .B2(n_1223), .ZN(n_894));
   XOR2_X1 i_855 (.A(n_1144), .B(n_1137), .Z(n_900));
   NAND2_X1 i_856 (.A1(n_1141), .A2(n_1138), .ZN(n_1137));
   NAND2_X1 i_857 (.A1(n_1143), .A2(n_1142), .ZN(n_1138));
   OR2_X1 i_858 (.A1(n_1143), .A2(n_1142), .ZN(n_1141));
   AOI21_X1 i_859 (.A(n_1270), .B1(n_1347), .B2(n_1266), .ZN(n_1142));
   AOI21_X1 i_860 (.A(n_1260), .B1(n_1339), .B2(n_1258), .ZN(n_1143));
   NAND2_X1 i_861 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [10]), .ZN(n_1144));
   XOR2_X1 i_862 (.A(n_1151), .B(n_1145), .Z(n_851));
   NAND2_X1 i_874 (.A1(n_1149), .A2(n_1148), .ZN(n_1145));
   NAND4_X1 i_875 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [9]), .A4(\r_weights[0] [1]), .ZN(n_1148));
   INV_X1 i_876 (.A(n_1150), .ZN(n_1149));
   AOI22_X1 i_877 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [9]), .B2(\r_weights[0] [1]), .ZN(n_1150));
   NAND2_X1 i_878 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [0]), .ZN(n_1151));
   XOR2_X1 i_879 (.A(n_1158), .B(n_1152), .Z(n_858));
   NAND2_X1 i_880 (.A1(n_1156), .A2(n_1155), .ZN(n_1152));
   NAND4_X1 i_881 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [6]), .A4(\r_weights[0] [4]), .ZN(n_1155));
   INV_X1 i_882 (.A(n_1157), .ZN(n_1156));
   AOI22_X1 i_883 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [6]), .B2(\r_weights[0] [4]), .ZN(n_1157));
   NAND2_X1 i_884 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [3]), .ZN(n_1158));
   XOR2_X1 i_885 (.A(n_1165), .B(n_1159), .Z(n_865));
   NAND2_X1 i_886 (.A1(n_1163), .A2(n_1162), .ZN(n_1159));
   NAND4_X1 i_887 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [8]), .A3(
      \r_values[0] [3]), .A4(\r_weights[0] [7]), .ZN(n_1162));
   INV_X1 i_888 (.A(n_1164), .ZN(n_1163));
   AOI22_X1 i_889 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [3]), .B2(\r_weights[0] [7]), .ZN(n_1164));
   NAND2_X1 i_890 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [6]), .ZN(n_1165));
   XOR2_X1 i_891 (.A(n_1203), .B(n_1166), .Z(n_872));
   NAND2_X1 i_892 (.A1(n_1170), .A2(n_1169), .ZN(n_1166));
   NAND3_X1 i_893 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [0]), .A3(n_1172), 
      .ZN(n_1169));
   INV_X1 i_894 (.A(n_1171), .ZN(n_1170));
   AOI21_X1 i_895 (.A(n_1172), .B1(\r_values[1] [10]), .B2(\r_weights[1] [0]), 
      .ZN(n_1171));
   AND2_X1 i_896 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [10]), .ZN(n_1172));
   NAND2_X1 i_897 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [9]), .ZN(n_1203));
   XOR2_X1 i_898 (.A(n_1252), .B(n_1204), .Z(n_879));
   AOI21_X1 i_899 (.A(n_1210), .B1(n_1339), .B2(n_1208), .ZN(n_1204));
   NAND2_X1 i_900 (.A1(n_1339), .A2(n_1208), .ZN(n_1207));
   INV_X1 i_901 (.A(n_1209), .ZN(n_1208));
   NAND2_X1 i_902 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [3]), .ZN(n_1209));
   AOI22_X1 i_903 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [3]), .B1(
      \r_values[1] [8]), .B2(\r_weights[1] [2]), .ZN(n_1210));
   XOR2_X1 i_904 (.A(n_1263), .B(n_1211), .Z(n_886));
   AOI21_X1 i_905 (.A(n_1217), .B1(n_1347), .B2(n_1215), .ZN(n_1211));
   NAND2_X1 i_906 (.A1(n_1347), .A2(n_1215), .ZN(n_1214));
   INV_X1 i_907 (.A(n_1216), .ZN(n_1215));
   NAND2_X1 i_908 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [6]), .ZN(n_1216));
   AOI22_X1 i_909 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [6]), .B1(
      \r_values[1] [5]), .B2(\r_weights[1] [5]), .ZN(n_1217));
   XOR2_X1 i_910 (.A(n_1271), .B(n_1218), .Z(n_893));
   AOI21_X1 i_911 (.A(n_1223), .B1(n_1353), .B2(n_1221), .ZN(n_1218));
   INV_X1 i_912 (.A(n_1222), .ZN(n_1221));
   NAND2_X1 i_913 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [9]), .ZN(n_1222));
   AOI22_X1 i_914 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [9]), .B1(
      \r_values[1] [2]), .B2(\r_weights[1] [8]), .ZN(n_1223));
   INV_X1 i_915 (.A(n_1224), .ZN(n_823));
   AOI22_X1 i_916 (.A1(n_1353), .A2(n_1312), .B1(n_1311), .B2(n_1307), .ZN(
      n_1224));
   OAI21_X1 i_917 (.A(n_1228), .B1(n_1231), .B2(n_1230), .ZN(n_782));
   OAI21_X1 i_918 (.A(n_1235), .B1(n_1238), .B2(n_1237), .ZN(n_789));
   OAI21_X1 i_919 (.A(n_1242), .B1(n_1245), .B2(n_1244), .ZN(n_796));
   AOI21_X1 i_920 (.A(n_1250), .B1(n_1256), .B2(n_1251), .ZN(n_803));
   XOR2_X1 i_921 (.A(n_1231), .B(n_1225), .Z(n_781));
   NAND2_X1 i_922 (.A1(n_1229), .A2(n_1228), .ZN(n_1225));
   NAND4_X1 i_923 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [8]), .A4(\r_weights[0] [1]), .ZN(n_1228));
   INV_X1 i_924 (.A(n_1230), .ZN(n_1229));
   AOI22_X1 i_925 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [8]), .B2(\r_weights[0] [1]), .ZN(n_1230));
   NAND2_X1 i_926 (.A1(\r_values[0] [9]), .A2(\r_weights[0] [0]), .ZN(n_1231));
   XOR2_X1 i_927 (.A(n_1238), .B(n_1232), .Z(n_788));
   NAND2_X1 i_928 (.A1(n_1236), .A2(n_1235), .ZN(n_1232));
   NAND4_X1 i_929 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [5]), .A4(\r_weights[0] [4]), .ZN(n_1235));
   INV_X1 i_943 (.A(n_1237), .ZN(n_1236));
   AOI22_X1 i_944 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [5]), .B2(\r_weights[0] [4]), .ZN(n_1237));
   NAND2_X1 i_945 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [3]), .ZN(n_1238));
   XOR2_X1 i_946 (.A(n_1245), .B(n_1239), .Z(n_795));
   NAND2_X1 i_947 (.A1(n_1243), .A2(n_1242), .ZN(n_1239));
   NAND3_X1 i_948 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [7]), .A3(n_1329), 
      .ZN(n_1242));
   INV_X1 i_949 (.A(n_1244), .ZN(n_1243));
   AOI21_X1 i_950 (.A(n_1329), .B1(\r_values[0] [2]), .B2(\r_weights[0] [7]), 
      .ZN(n_1244));
   NAND2_X1 i_951 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [6]), .ZN(n_1245));
   XOR2_X1 i_952 (.A(n_1256), .B(n_1246), .Z(n_802));
   NAND2_X1 i_953 (.A1(n_1251), .A2(n_1249), .ZN(n_1246));
   INV_X1 i_954 (.A(n_1250), .ZN(n_1249));
   AOI22_X1 i_955 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [1]), .B1(
      \r_values[1] [9]), .B2(\r_weights[1] [0]), .ZN(n_1250));
   NAND2_X1 i_956 (.A1(n_1341), .A2(n_1252), .ZN(n_1251));
   INV_X1 i_957 (.A(n_1253), .ZN(n_1252));
   NAND2_X1 i_958 (.A1(\r_values[1] [9]), .A2(\r_weights[1] [1]), .ZN(n_1253));
   NAND2_X1 i_959 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [9]), .ZN(n_1256));
   XOR2_X1 i_960 (.A(n_1339), .B(n_1257), .Z(n_809));
   NOR2_X1 i_961 (.A1(n_1260), .A2(n_1259), .ZN(n_1257));
   INV_X1 i_962 (.A(n_1259), .ZN(n_1258));
   AOI22_X1 i_963 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [4]), .B1(
      \r_values[1] [6]), .B2(\r_weights[1] [3]), .ZN(n_1259));
   NOR2_X1 i_964 (.A1(n_1428), .A2(n_1264), .ZN(n_1260));
   INV_X1 i_965 (.A(n_1264), .ZN(n_1263));
   NAND2_X1 i_966 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [4]), .ZN(n_1264));
   XOR2_X1 i_967 (.A(n_1347), .B(n_1265), .Z(n_816));
   NOR2_X1 i_968 (.A1(n_1270), .A2(n_1267), .ZN(n_1265));
   INV_X1 i_969 (.A(n_1267), .ZN(n_1266));
   AOI22_X1 i_970 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [7]), .B1(
      \r_values[1] [3]), .B2(\r_weights[1] [6]), .ZN(n_1267));
   AND2_X1 i_971 (.A1(n_1434), .A2(n_1271), .ZN(n_1270));
   INV_X1 i_972 (.A(n_1272), .ZN(n_1271));
   NAND2_X1 i_973 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [7]), .ZN(n_1272));
   XOR2_X1 i_974 (.A(n_1311), .B(n_1307), .Z(n_822));
   NOR2_X1 i_975 (.A1(n_1355), .A2(n_1308), .ZN(n_1307));
   NOR2_X1 i_976 (.A1(n_1434), .A2(n_1350), .ZN(n_1308));
   XNOR2_X1 i_977 (.A(n_1354), .B(n_1312), .ZN(n_1311));
   AND2_X1 i_978 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [9]), .ZN(n_1312));
   OAI21_X1 i_979 (.A(n_1314), .B1(n_1319), .B2(n_1318), .ZN(n_722));
   OAI21_X1 i_980 (.A(n_1321), .B1(n_1326), .B2(n_1325), .ZN(n_729));
   OAI21_X1 i_981 (.A(n_1328), .B1(n_1334), .B2(n_1333), .ZN(n_736));
   OAI21_X1 i_982 (.A(n_1336), .B1(n_1342), .B2(n_1340), .ZN(n_743));
   OAI21_X1 i_983 (.A(n_1346), .B1(n_1428), .B2(n_1348), .ZN(n_750));
   XOR2_X1 i_984 (.A(n_1319), .B(n_1313), .Z(n_721));
   NAND2_X1 i_985 (.A1(n_1315), .A2(n_1314), .ZN(n_1313));
   NAND4_X1 i_986 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [7]), .A4(\r_weights[0] [1]), .ZN(n_1314));
   INV_X1 i_987 (.A(n_1318), .ZN(n_1315));
   AOI22_X1 i_988 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [7]), .B2(\r_weights[0] [1]), .ZN(n_1318));
   NAND2_X1 i_989 (.A1(\r_values[0] [8]), .A2(\r_weights[0] [0]), .ZN(n_1319));
   XOR2_X1 i_990 (.A(n_1326), .B(n_1320), .Z(n_728));
   NAND2_X1 i_991 (.A1(n_1322), .A2(n_1321), .ZN(n_1320));
   NAND4_X1 i_992 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [4]), .A4(\r_weights[0] [4]), .ZN(n_1321));
   INV_X1 i_993 (.A(n_1325), .ZN(n_1322));
   AOI22_X1 i_994 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [4]), .ZN(n_1325));
   NAND2_X1 i_995 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [3]), .ZN(n_1326));
   XOR2_X1 i_996 (.A(n_1334), .B(n_1327), .Z(n_735));
   NAND2_X1 i_997 (.A1(n_1332), .A2(n_1328), .ZN(n_1327));
   NAND2_X1 i_998 (.A1(n_1421), .A2(n_1329), .ZN(n_1328));
   AND2_X1 i_999 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [8]), .ZN(n_1329));
   INV_X1 i_1000 (.A(n_1333), .ZN(n_1332));
   AOI22_X1 i_1001 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [8]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [7]), .ZN(n_1333));
   NAND2_X1 i_1002 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [6]), .ZN(n_1334));
   XOR2_X1 i_1003 (.A(n_1341), .B(n_1335), .Z(n_742));
   AOI21_X1 i_1004 (.A(n_1340), .B1(n_1457), .B2(n_1339), .ZN(n_1335));
   NAND2_X1 i_1005 (.A1(n_1457), .A2(n_1339), .ZN(n_1336));
   AND2_X1 i_1006 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [2]), .ZN(n_1339));
   AOI22_X1 i_1021 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [2]), .B1(
      \r_values[1] [7]), .B2(\r_weights[1] [1]), .ZN(n_1340));
   INV_X1 i_1022 (.A(n_1342), .ZN(n_1341));
   NAND2_X1 i_1023 (.A1(\r_values[1] [8]), .A2(\r_weights[1] [0]), .ZN(n_1342));
   XOR2_X1 i_1024 (.A(n_1427), .B(n_1343), .Z(n_749));
   AOI21_X1 i_1025 (.A(n_1348), .B1(n_1467), .B2(n_1347), .ZN(n_1343));
   NAND2_X1 i_1026 (.A1(n_1467), .A2(n_1347), .ZN(n_1346));
   AND2_X1 i_1027 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [5]), .ZN(n_1347));
   AOI22_X1 i_1028 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [5]), .B1(
      \r_values[1] [4]), .B2(\r_weights[1] [4]), .ZN(n_1348));
   XOR2_X1 i_1029 (.A(n_1434), .B(n_1349), .Z(n_756));
   NOR2_X1 i_1030 (.A1(n_1355), .A2(n_1350), .ZN(n_1349));
   NOR2_X1 i_1031 (.A1(n_1364), .A2(n_1354), .ZN(n_1350));
   INV_X1 i_1032 (.A(n_1354), .ZN(n_1353));
   NAND2_X1 i_1033 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [8]), .ZN(n_1354));
   AOI22_X1 i_1034 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [8]), .B1(
      \r_values[1] [1]), .B2(\r_weights[1] [7]), .ZN(n_1355));
   AOI21_X1 i_1035 (.A(n_1360), .B1(n_1364), .B2(n_1357), .ZN(n_700));
   OAI21_X1 i_1036 (.A(n_1368), .B1(n_1371), .B2(n_1370), .ZN(n_665));
   OAI21_X1 i_1037 (.A(n_1375), .B1(n_1380), .B2(n_1377), .ZN(n_672));
   AOI21_X1 i_1038 (.A(n_1384), .B1(n_1422), .B2(n_1382), .ZN(n_679));
   OAI21_X1 i_1039 (.A(n_1426), .B1(n_1460), .B2(n_1429), .ZN(n_686));
   OAI21_X1 i_1040 (.A(n_1433), .B1(n_1468), .B2(n_1435), .ZN(n_693));
   XOR2_X1 i_1041 (.A(n_1364), .B(n_1356), .Z(n_699));
   OAI21_X1 i_1042 (.A(n_1357), .B1(n_1363), .B2(n_1361), .ZN(n_1356));
   NAND2_X1 i_1043 (.A1(n_1363), .A2(n_1361), .ZN(n_1357));
   NOR2_X1 i_1044 (.A1(n_1363), .A2(n_1361), .ZN(n_1360));
   NOR2_X1 i_1045 (.A1(n_1463), .A2(n_1362), .ZN(n_1361));
   NOR2_X1 i_1046 (.A1(n_1529), .A2(n_1464), .ZN(n_1362));
   AOI21_X1 i_1047 (.A(n_1455), .B1(n_1461), .B2(n_1456), .ZN(n_1363));
   NAND2_X1 i_1048 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [7]), .ZN(n_1364));
   XOR2_X1 i_1049 (.A(n_1371), .B(n_1367), .Z(n_664));
   NAND2_X1 i_1050 (.A1(n_1369), .A2(n_1368), .ZN(n_1367));
   NAND4_X1 i_1051 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [6]), .A4(\r_weights[0] [1]), .ZN(n_1368));
   INV_X1 i_1052 (.A(n_1370), .ZN(n_1369));
   AOI22_X1 i_1053 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [6]), .B2(\r_weights[0] [1]), .ZN(n_1370));
   NAND2_X1 i_1054 (.A1(\r_values[0] [7]), .A2(\r_weights[0] [0]), .ZN(n_1371));
   XOR2_X1 i_1055 (.A(n_1380), .B(n_1374), .Z(n_671));
   NAND2_X1 i_1056 (.A1(n_1376), .A2(n_1375), .ZN(n_1374));
   NAND4_X1 i_1057 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [5]), .A3(
      \r_values[0] [3]), .A4(\r_weights[0] [4]), .ZN(n_1375));
   INV_X1 i_1058 (.A(n_1377), .ZN(n_1376));
   AOI22_X1 i_1059 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [3]), .B2(\r_weights[0] [4]), .ZN(n_1377));
   NAND2_X1 i_1060 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [3]), .ZN(n_1380));
   XOR2_X1 i_1061 (.A(n_1422), .B(n_1381), .Z(n_678));
   NAND2_X1 i_1062 (.A1(n_1383), .A2(n_1382), .ZN(n_1381));
   NAND3_X1 i_1063 (.A1(\r_values[1] [7]), .A2(\r_weights[1] [0]), .A3(n_1421), 
      .ZN(n_1382));
   INV_X1 i_1064 (.A(n_1384), .ZN(n_1383));
   AOI21_X1 i_1065 (.A(n_1421), .B1(\r_values[1] [7]), .B2(\r_weights[1] [0]), 
      .ZN(n_1384));
   AND2_X1 i_1066 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [7]), .ZN(n_1421));
   NAND2_X1 i_1067 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [6]), .ZN(n_1422));
   XOR2_X1 i_1068 (.A(n_1457), .B(n_1425), .Z(n_685));
   AOI21_X1 i_1069 (.A(n_1429), .B1(n_1529), .B2(n_1427), .ZN(n_1425));
   NAND2_X1 i_1070 (.A1(n_1529), .A2(n_1427), .ZN(n_1426));
   INV_X1 i_1071 (.A(n_1428), .ZN(n_1427));
   NAND2_X1 i_1072 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [3]), .ZN(n_1428));
   AOI22_X1 i_1073 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [3]), .B1(
      \r_values[1] [5]), .B2(\r_weights[1] [2]), .ZN(n_1429));
   XOR2_X1 i_1074 (.A(n_1467), .B(n_1432), .Z(n_692));
   AOI21_X1 i_1075 (.A(n_1435), .B1(n_1537), .B2(n_1434), .ZN(n_1432));
   NAND2_X1 i_1076 (.A1(n_1537), .A2(n_1434), .ZN(n_1433));
   AND2_X1 i_1077 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [6]), .ZN(n_1434));
   AOI22_X1 i_1078 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [6]), .B1(
      \r_values[1] [2]), .B2(\r_weights[1] [5]), .ZN(n_1435));
   INV_X1 i_1079 (.A(n_1436), .ZN(n_644));
   AOI22_X1 i_1080 (.A1(n_1537), .A2(n_1474), .B1(n_1471), .B2(n_1469), .ZN(
      n_1436));
   OAI21_X1 i_1081 (.A(n_1440), .B1(n_1443), .B2(n_1442), .ZN(n_617));
   OAI21_X1 i_1082 (.A(n_1447), .B1(n_1450), .B2(n_1449), .ZN(n_624));
   XOR2_X1 i_1083 (.A(n_1443), .B(n_1439), .Z(n_616));
   NAND2_X1 i_1084 (.A1(n_1441), .A2(n_1440), .ZN(n_1439));
   NAND4_X1 i_1085 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [5]), .A4(\r_weights[0] [1]), .ZN(n_1440));
   INV_X1 i_1086 (.A(n_1442), .ZN(n_1441));
   AOI22_X1 i_1087 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [5]), .B2(\r_weights[0] [1]), .ZN(n_1442));
   NAND2_X1 i_1088 (.A1(\r_values[0] [6]), .A2(\r_weights[0] [0]), .ZN(n_1443));
   XOR2_X1 i_1089 (.A(n_1450), .B(n_1446), .Z(n_623));
   NAND2_X1 i_1090 (.A1(n_1448), .A2(n_1447), .ZN(n_1446));
   NAND3_X1 i_1091 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [4]), .A3(n_1484), 
      .ZN(n_1447));
   INV_X1 i_1107 (.A(n_1449), .ZN(n_1448));
   AOI21_X1 i_1108 (.A(n_1484), .B1(\r_values[0] [2]), .B2(\r_weights[0] [4]), 
      .ZN(n_1449));
   NAND2_X1 i_1109 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [3]), .ZN(n_1450));
   XOR2_X1 i_1110 (.A(n_1461), .B(n_1453), .Z(n_630));
   NAND2_X1 i_1111 (.A1(n_1456), .A2(n_1454), .ZN(n_1453));
   INV_X1 i_1112 (.A(n_1455), .ZN(n_1454));
   AOI22_X1 i_1113 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [1]), .B1(
      \r_values[1] [6]), .B2(\r_weights[1] [0]), .ZN(n_1455));
   NAND2_X1 i_1114 (.A1(n_1533), .A2(n_1457), .ZN(n_1456));
   INV_X1 i_1115 (.A(n_1460), .ZN(n_1457));
   NAND2_X1 i_1116 (.A1(\r_values[1] [6]), .A2(\r_weights[1] [1]), .ZN(n_1460));
   NAND2_X1 i_1117 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [6]), .ZN(n_1461));
   XOR2_X1 i_1118 (.A(n_1529), .B(n_1462), .Z(n_637));
   NOR2_X1 i_1119 (.A1(n_1464), .A2(n_1463), .ZN(n_1462));
   AOI22_X1 i_1120 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [4]), .B1(
      \r_values[1] [3]), .B2(\r_weights[1] [3]), .ZN(n_1463));
   AND2_X1 i_1121 (.A1(n_1569), .A2(n_1467), .ZN(n_1464));
   INV_X1 i_1122 (.A(n_1468), .ZN(n_1467));
   NAND2_X1 i_1123 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [4]), .ZN(n_1468));
   XOR2_X1 i_1124 (.A(n_1471), .B(n_1469), .Z(n_643));
   NOR2_X1 i_1125 (.A1(n_1541), .A2(n_1470), .ZN(n_1469));
   NOR2_X1 i_1126 (.A1(n_1569), .A2(n_1536), .ZN(n_1470));
   XNOR2_X1 i_1127 (.A(n_1540), .B(n_1474), .ZN(n_1471));
   AND2_X1 i_1128 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [6]), .ZN(n_1474));
   OAI21_X1 i_1129 (.A(n_1476), .B1(n_1481), .B2(n_1478), .ZN(n_579));
   OAI21_X1 i_1130 (.A(n_1483), .B1(n_1488), .B2(n_1487), .ZN(n_586));
   OAI21_X1 i_1131 (.A(n_1490), .B1(n_1534), .B2(n_1530), .ZN(n_593));
   XOR2_X1 i_1132 (.A(n_1481), .B(n_1475), .Z(n_578));
   NAND2_X1 i_1133 (.A1(n_1477), .A2(n_1476), .ZN(n_1475));
   NAND4_X1 i_1134 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [4]), .A4(\r_weights[0] [1]), .ZN(n_1476));
   INV_X1 i_1135 (.A(n_1478), .ZN(n_1477));
   AOI22_X1 i_1136 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [4]), .B2(\r_weights[0] [1]), .ZN(n_1478));
   NAND2_X1 i_1137 (.A1(\r_values[0] [5]), .A2(\r_weights[0] [0]), .ZN(n_1481));
   XOR2_X1 i_1138 (.A(n_1488), .B(n_1482), .Z(n_585));
   NAND2_X1 i_1139 (.A1(n_1485), .A2(n_1483), .ZN(n_1482));
   NAND2_X1 i_1140 (.A1(n_1563), .A2(n_1484), .ZN(n_1483));
   AND2_X1 i_1141 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [5]), .ZN(n_1484));
   INV_X1 i_1142 (.A(n_1487), .ZN(n_1485));
   AOI22_X1 i_1143 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [5]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [4]), .ZN(n_1487));
   NAND2_X1 i_1144 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [3]), .ZN(n_1488));
   XOR2_X1 i_1145 (.A(n_1533), .B(n_1489), .Z(n_592));
   AOI21_X1 i_1146 (.A(n_1530), .B1(n_1585), .B2(n_1529), .ZN(n_1489));
   NAND2_X1 i_1147 (.A1(n_1585), .A2(n_1529), .ZN(n_1490));
   AND2_X1 i_1148 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [2]), .ZN(n_1529));
   AOI22_X1 i_1149 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [2]), .B1(
      \r_values[1] [4]), .B2(\r_weights[1] [1]), .ZN(n_1530));
   INV_X1 i_1150 (.A(n_1534), .ZN(n_1533));
   NAND2_X1 i_1151 (.A1(\r_values[1] [5]), .A2(\r_weights[1] [0]), .ZN(n_1534));
   XOR2_X1 i_1152 (.A(n_1569), .B(n_1535), .Z(n_599));
   NOR2_X1 i_1153 (.A1(n_1541), .A2(n_1536), .ZN(n_1535));
   NOR2_X1 i_1154 (.A1(n_1549), .A2(n_1540), .ZN(n_1536));
   INV_X1 i_1155 (.A(n_1540), .ZN(n_1537));
   NAND2_X1 i_1156 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [5]), .ZN(n_1540));
   AOI22_X1 i_1157 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [5]), .B1(
      \r_values[1] [1]), .B2(\r_weights[1] [4]), .ZN(n_1541));
   AOI21_X1 i_1158 (.A(n_1544), .B1(n_1549), .B2(n_1543), .ZN(n_565));
   OAI21_X1 i_1159 (.A(n_1551), .B1(n_1556), .B2(n_1555), .ZN(n_544));
   AOI21_X1 i_1160 (.A(n_1562), .B1(n_1564), .B2(n_1558), .ZN(n_551));
   OAI21_X1 i_1161 (.A(n_1568), .B1(n_1586), .B2(n_1570), .ZN(n_558));
   XOR2_X1 i_1162 (.A(n_1549), .B(n_1542), .Z(n_564));
   OAI21_X1 i_1163 (.A(n_1543), .B1(n_1548), .B2(n_1547), .ZN(n_1542));
   NAND2_X1 i_1164 (.A1(n_1548), .A2(n_1547), .ZN(n_1543));
   NOR2_X1 i_1165 (.A1(n_1548), .A2(n_1547), .ZN(n_1544));
   OAI21_X1 i_1166 (.A(n_1575), .B1(n_1578), .B2(n_1577), .ZN(n_1547));
   AOI21_X1 i_1167 (.A(n_1583), .B1(n_1589), .B2(n_1584), .ZN(n_1548));
   NAND2_X1 i_1168 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [4]), .ZN(n_1549));
   XOR2_X1 i_1169 (.A(n_1556), .B(n_1550), .Z(n_543));
   NAND2_X1 i_1170 (.A1(n_1554), .A2(n_1551), .ZN(n_1550));
   NAND4_X1 i_1171 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [3]), .A4(\r_weights[0] [1]), .ZN(n_1551));
   INV_X1 i_1172 (.A(n_1555), .ZN(n_1554));
   AOI22_X1 i_1173 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [3]), .B2(\r_weights[0] [1]), .ZN(n_1555));
   NAND2_X1 i_1174 (.A1(\r_values[0] [4]), .A2(\r_weights[0] [0]), .ZN(n_1556));
   XOR2_X1 i_1175 (.A(n_1564), .B(n_1557), .Z(n_550));
   NAND2_X1 i_1176 (.A1(n_1561), .A2(n_1558), .ZN(n_1557));
   NAND3_X1 i_1194 (.A1(\r_values[1] [4]), .A2(\r_weights[1] [0]), .A3(n_1563), 
      .ZN(n_1558));
   INV_X1 i_1195 (.A(n_1562), .ZN(n_1561));
   AOI21_X1 i_1196 (.A(n_1563), .B1(\r_values[1] [4]), .B2(\r_weights[1] [0]), 
      .ZN(n_1562));
   AND2_X1 i_1197 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [4]), .ZN(n_1563));
   NAND2_X1 i_1198 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [3]), .ZN(n_1564));
   XOR2_X1 i_1199 (.A(n_1585), .B(n_1565), .Z(n_557));
   AOI21_X1 i_1200 (.A(n_1570), .B1(n_1640), .B2(n_1569), .ZN(n_1565));
   NAND2_X1 i_1201 (.A1(n_1640), .A2(n_1569), .ZN(n_1568));
   AND2_X1 i_1202 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [3]), .ZN(n_1569));
   AOI22_X1 i_1203 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [3]), .B1(
      \r_values[1] [2]), .B2(\r_weights[1] [2]), .ZN(n_1570));
   INV_X1 i_1204 (.A(n_1571), .ZN(n_531));
   AOI22_X1 i_1205 (.A1(n_1640), .A2(n_1592), .B1(n_1591), .B2(n_1590), .ZN(
      n_1571));
   XOR2_X1 i_1206 (.A(n_1578), .B(n_1572), .Z(n_517));
   NAND2_X1 i_1207 (.A1(n_1576), .A2(n_1575), .ZN(n_1572));
   NAND4_X1 i_1208 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [2]), .A4(\r_weights[0] [1]), .ZN(n_1575));
   INV_X1 i_1209 (.A(n_1577), .ZN(n_1576));
   AOI22_X1 i_1210 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [2]), .B2(\r_weights[0] [1]), .ZN(n_1577));
   NAND2_X1 i_1211 (.A1(\r_values[0] [3]), .A2(\r_weights[0] [0]), .ZN(n_1578));
   XOR2_X1 i_1212 (.A(n_1589), .B(n_1579), .Z(n_524));
   NAND2_X1 i_1213 (.A1(n_1584), .A2(n_1582), .ZN(n_1579));
   INV_X1 i_1214 (.A(n_1583), .ZN(n_1582));
   AOI22_X1 i_1215 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [1]), .B1(
      \r_values[1] [3]), .B2(\r_weights[1] [0]), .ZN(n_1583));
   NAND2_X1 i_1216 (.A1(n_1643), .A2(n_1585), .ZN(n_1584));
   INV_X1 i_1217 (.A(n_1586), .ZN(n_1585));
   NAND2_X1 i_1218 (.A1(\r_values[1] [3]), .A2(\r_weights[1] [1]), .ZN(n_1586));
   NAND2_X1 i_1219 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [3]), .ZN(n_1589));
   XOR2_X1 i_1220 (.A(n_1591), .B(n_1590), .Z(n_530));
   OAI21_X1 i_1221 (.A(n_1637), .B1(n_1644), .B2(n_1642), .ZN(n_1590));
   XNOR2_X1 i_1222 (.A(n_1641), .B(n_1592), .ZN(n_1591));
   AND2_X1 i_1223 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [3]), .ZN(n_1592));
   OAI21_X1 i_1224 (.A(n_1596), .B1(n_1598), .B2(n_1593), .ZN(n_502));
   NAND2_X1 i_1225 (.A1(\r_values[0] [2]), .A2(\r_weights[0] [0]), .ZN(n_1593));
   NAND4_X1 i_1226 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [2]), .A3(
      \r_values[0] [1]), .A4(\r_weights[0] [1]), .ZN(n_1596));
   INV_X1 i_1227 (.A(n_1598), .ZN(n_1597));
   AOI22_X1 i_1228 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [2]), .B1(
      \r_values[0] [1]), .B2(\r_weights[0] [1]), .ZN(n_1598));
   XOR2_X1 i_1229 (.A(n_1643), .B(n_1599), .Z(n_508));
   NOR2_X1 i_1230 (.A1(n_1642), .A2(n_1636), .ZN(n_1599));
   INV_X1 i_1231 (.A(n_1637), .ZN(n_1636));
   NAND3_X1 i_1232 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [1]), .A3(n_1640), 
      .ZN(n_1637));
   INV_X1 i_1233 (.A(n_1641), .ZN(n_1640));
   NAND2_X1 i_1234 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [2]), .ZN(n_1641));
   AOI22_X1 i_1235 (.A1(\r_values[1] [0]), .A2(\r_weights[1] [2]), .B1(
      \r_values[1] [1]), .B2(\r_weights[1] [1]), .ZN(n_1642));
   INV_X1 i_1236 (.A(n_1644), .ZN(n_1643));
   NAND2_X1 i_1237 (.A1(\r_values[1] [2]), .A2(\r_weights[1] [0]), .ZN(n_1644));
   OAI22_X1 i_1238 (.A1(n_1650), .A2(n_1649), .B1(n_1648), .B2(n_1647), .ZN(
      n_495));
   XNOR2_X1 i_1239 (.A(n_1650), .B(n_1649), .ZN(n_1647));
   NAND2_X1 i_1240 (.A1(\r_values[0] [1]), .A2(\r_weights[0] [0]), .ZN(n_1648));
   NAND2_X1 i_1241 (.A1(\r_values[1] [1]), .A2(\r_weights[1] [0]), .ZN(n_1649));
   NAND2_X1 i_1242 (.A1(\r_values[0] [0]), .A2(\r_weights[0] [1]), .ZN(n_1650));
   XOR2_X1 i_1243 (.A(n_1695), .B(n_1651), .Z(\sums[2] [26]));
   XNOR2_X1 i_1244 (.A(n_1675), .B(n_1654), .ZN(n_1651));
   XNOR2_X1 i_1245 (.A(n_1665), .B(n_1655), .ZN(n_1654));
   AOI21_X1 i_1246 (.A(n_1661), .B1(n_1662), .B2(n_1657), .ZN(n_1655));
   INV_X1 i_1247 (.A(n_1657), .ZN(n_1656));
   NAND2_X1 i_1248 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [10]), .ZN(n_1657));
   INV_X1 i_1249 (.A(n_1661), .ZN(n_1658));
   AOI22_X1 i_1250 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [12]), .B1(
      \r_values[1] [14]), .B2(\r_weights[1] [11]), .ZN(n_1661));
   OR2_X1 i_1251 (.A1(n_1758), .A2(n_1664), .ZN(n_1662));
   INV_X1 i_1252 (.A(n_1664), .ZN(n_1663));
   NAND2_X1 i_1253 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [11]), .ZN(n_1664));
   AOI21_X1 i_1254 (.A(n_1670), .B1(n_1671), .B2(n_1668), .ZN(n_1665));
   NAND2_X1 i_1255 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [10]), .ZN(n_1668));
   INV_X1 i_1256 (.A(n_1670), .ZN(n_1669));
   AOI22_X1 i_1257 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [12]), .B1(
      \r_values[0] [14]), .B2(\r_weights[0] [11]), .ZN(n_1670));
   NAND3_X1 i_1258 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [12]), .A3(n_1672), 
      .ZN(n_1671));
   AND2_X1 i_1259 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [11]), .ZN(n_1672));
   XNOR2_X1 i_1260 (.A(n_1684), .B(n_1676), .ZN(n_1675));
   AOI21_X1 i_1261 (.A(n_1679), .B1(n_1682), .B2(n_1677), .ZN(n_1676));
   NAND2_X1 i_1262 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [13]), .ZN(n_1677));
   INV_X1 i_1263 (.A(n_1679), .ZN(n_1678));
   AOI22_X1 i_1264 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [15]), .B1(
      \r_values[0] [11]), .B2(\r_weights[0] [14]), .ZN(n_1679));
   NAND3_X1 i_1265 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [15]), .A3(n_1683), 
      .ZN(n_1682));
   AND2_X1 i_1266 (.A1(\r_values[0] [10]), .A2(\r_weights[0] [14]), .ZN(n_1683));
   AOI21_X1 i_1267 (.A(n_1690), .B1(n_1691), .B2(n_1686), .ZN(n_1684));
   INV_X1 i_1268 (.A(n_1686), .ZN(n_1685));
   NAND2_X1 i_1269 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [13]), .ZN(n_1686));
   INV_X1 i_1270 (.A(n_1690), .ZN(n_1689));
   AOI22_X1 i_1271 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [15]), .B1(
      \r_values[1] [11]), .B2(\r_weights[1] [14]), .ZN(n_1690));
   NAND3_X1 i_1290 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [15]), .A3(n_1692), 
      .ZN(n_1691));
   AND2_X1 i_1291 (.A1(\r_values[1] [10]), .A2(\r_weights[1] [14]), .ZN(n_1692));
   XNOR2_X1 i_1292 (.A(n_1697), .B(n_1696), .ZN(n_1695));
   XNOR2_X1 i_1293 (.A(n_1751), .B(n_1698), .ZN(n_1696));
   XOR2_X1 i_1294 (.A(n_1762), .B(n_1743), .Z(n_1697));
   XNOR2_X1 i_1295 (.A(n_1740), .B(n_1699), .ZN(n_1698));
   XOR2_X1 i_1296 (.A(n_1737), .B(n_1736), .Z(n_1699));
   NAND2_X1 i_1297 (.A1(\r_values[0] [14]), .A2(\r_weights[0] [12]), .ZN(n_1736));
   NAND2_X1 i_1298 (.A1(\r_values[1] [12]), .A2(\r_weights[1] [14]), .ZN(n_1737));
   XNOR2_X1 i_1299 (.A(n_1742), .B(n_1741), .ZN(n_1740));
   NAND2_X1 i_1300 (.A1(\r_values[0] [11]), .A2(\r_weights[0] [15]), .ZN(n_1741));
   AND2_X1 i_1301 (.A1(\r_values[1] [13]), .A2(\r_weights[1] [13]), .ZN(n_1742));
   XOR2_X1 i_1302 (.A(n_1748), .B(n_1744), .Z(n_1743));
   XNOR2_X1 i_1303 (.A(n_173), .B(n_1747), .ZN(n_1744));
   XNOR2_X1 i_1304 (.A(\sums[0] [26]), .B(n_169), .ZN(n_1747));
   XNOR2_X1 i_1305 (.A(n_1750), .B(n_1749), .ZN(n_1748));
   XNOR2_X1 i_1306 (.A(n_175), .B(n_177), .ZN(n_1749));
   AND2_X1 i_1307 (.A1(\r_values[0] [13]), .A2(\r_weights[0] [13]), .ZN(n_1750));
   XOR2_X1 i_1308 (.A(n_1757), .B(n_1754), .Z(n_1751));
   XNOR2_X1 i_1309 (.A(n_1756), .B(n_1755), .ZN(n_1754));
   NAND2_X1 i_1310 (.A1(\r_values[0] [15]), .A2(\r_weights[0] [11]), .ZN(n_1755));
   NAND2_X1 i_1311 (.A1(\r_values[1] [11]), .A2(\r_weights[1] [15]), .ZN(n_1756));
   XNOR2_X1 i_1312 (.A(n_1761), .B(n_1758), .ZN(n_1757));
   NAND2_X1 i_1313 (.A1(\r_values[1] [14]), .A2(\r_weights[1] [12]), .ZN(n_1758));
   AND2_X1 i_1314 (.A1(\r_values[1] [15]), .A2(\r_weights[1] [11]), .ZN(n_1761));
   XOR2_X1 i_1315 (.A(n_1768), .B(n_1763), .Z(n_1762));
   XNOR2_X1 i_1316 (.A(n_1765), .B(n_1764), .ZN(n_1763));
   XOR2_X1 i_1317 (.A(n_161), .B(n_163), .Z(n_1764));
   NAND2_X1 i_1318 (.A1(\r_values[0] [12]), .A2(\r_weights[0] [14]), .ZN(n_1765));
   XNOR2_X1 i_1319 (.A(n_1770), .B(n_1769), .ZN(n_1768));
   XOR2_X1 i_1320 (.A(n_165), .B(n_167), .Z(n_1769));
   XOR2_X1 i_1321 (.A(n_171), .B(n_210), .Z(n_1770));
   INV_X1 i_1322 (.A(\sums[0] [12]), .ZN(n_1771));
   INV_X1 i_1323 (.A(\sums[0] [13]), .ZN(n_1772));
   INV_X1 i_1324 (.A(\sums[0] [15]), .ZN(n_1775));
   INV_X1 i_1325 (.A(\sums[0] [18]), .ZN(n_1776));
   INV_X1 i_1326 (.A(\sums[0] [21]), .ZN(n_1777));
   INV_X1 i_1327 (.A(\sums[0] [24]), .ZN(n_1778));
endmodule

module ALU(clk, \i_values[0] , \i_values[1] , i_single, load_enable, clear, value);
   input clk;
   input [15:0]\i_values[0] ;
   input [15:0]\i_values[1] ;
   input [15:0]i_single;
   input [1:0]load_enable;
   input clear;
   output [15:0]value;

   wire [15:0]\r_values[0] ;
   wire [15:0]\r_values[1] ;
   wire [15:0]\r_weights[0] ;
   wire [15:0]\r_weights[1] ;
   wire [15:0]r_bias;
   wire n_0_0;
   wire n_0_1_0;
   wire n_0_1;
   wire n_0_1_1;
   wire n_0_2;
   wire n_0_1_2;
   wire n_0_3;
   wire n_0_1_3;
   wire n_0_4;
   wire n_0_1_4;
   wire n_0_5;
   wire n_0_1_5;
   wire n_0_6;
   wire n_0_1_6;
   wire n_0_7;
   wire n_0_1_7;
   wire n_0_8;
   wire n_0_1_8;
   wire n_0_9;
   wire n_0_1_9;
   wire n_0_10;
   wire n_0_1_10;
   wire n_0_11;
   wire n_0_1_11;
   wire n_0_12;
   wire n_0_1_12;
   wire n_0_13;
   wire n_0_1_13;
   wire n_0_14;
   wire n_0_1_14;
   wire n_0_15;
   wire n_0_1_15;
   wire n_0_16;
   wire n_0_1_16;
   wire n_0_17;
   wire n_0_1_17;
   wire n_0_18;
   wire n_0_1_18;
   wire n_0_19;
   wire n_0_1_19;
   wire n_0_20;
   wire n_0_1_20;
   wire n_0_21;
   wire n_0_1_21;
   wire n_0_22;
   wire n_0_1_22;
   wire n_0_23;
   wire n_0_1_23;
   wire n_0_24;
   wire n_0_1_24;
   wire n_0_25;
   wire n_0_1_25;
   wire n_0_26;
   wire n_0_1_26;
   wire n_0_27;
   wire n_0_1_27;
   wire n_0_28;
   wire n_0_1_28;
   wire n_0_29;
   wire n_0_1_29;
   wire n_0_30;
   wire n_0_1_30;
   wire n_0_31;
   wire n_0_1_31;
   wire n_0_32;
   wire n_0_1_32;
   wire n_0_33;
   wire n_0_1_33;
   wire n_0_34;
   wire n_0_1_34;
   wire n_0_35;
   wire n_0_1_35;
   wire n_0_36;
   wire n_0_1_36;
   wire n_0_37;
   wire n_0_1_37;
   wire n_0_38;
   wire n_0_1_38;
   wire n_0_39;
   wire n_0_1_39;
   wire n_0_40;
   wire n_0_1_40;
   wire n_0_41;
   wire n_0_1_41;
   wire n_0_42;
   wire n_0_1_42;
   wire n_0_43;
   wire n_0_1_43;
   wire n_0_44;
   wire n_0_1_44;
   wire n_0_45;
   wire n_0_1_45;
   wire n_0_46;
   wire n_0_1_46;
   wire n_0_47;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_48;
   wire n_0_49;
   wire n_0_80;
   wire n_0_79;
   wire n_0_78;
   wire n_0_77;
   wire n_0_76;
   wire n_0_75;
   wire n_0_74;
   wire n_0_73;
   wire n_0_71;
   wire n_0_70;
   wire n_0_69;
   wire n_0_68;
   wire n_0_67;
   wire n_0_66;
   wire n_0_65;
   wire n_0_64;
   wire n_0_63;
   wire n_0_62;
   wire n_0_61;
   wire n_0_60;
   wire n_0_59;
   wire n_0_58;
   wire n_0_57;
   wire n_0_56;
   wire n_0_55;
   wire n_0_54;
   wire n_0_53;
   wire n_0_52;
   wire n_0_51;
   wire n_0_50;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_1_52;
   wire n_0_72;

   datapath i_0_0 (.\sums[0] ({r_bias[15], r_bias[14], r_bias[13], r_bias[12], 
      r_bias[11], r_bias[10], r_bias[9], r_bias[8], r_bias[7], r_bias[6], 
      r_bias[5], r_bias[4], r_bias[3], r_bias[2], r_bias[1], r_bias[0], 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .\sums[2] ({
      value[15], value[14], value[13], value[12], value[11], value[10], value[9], 
      value[8], value[7], value[6], value[5], value[4], value[3], value[2], 
      value[1], value[0], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10}), .\r_values[0] (\r_values[0] ), .\r_weights[0] (
      \r_weights[0] ), .\r_values[1] (\r_values[1] ), .\r_weights[1] (
      \r_weights[1] ));
   DFF_X1 \r_values_reg[0][15]  (.D(n_0_50), .CK(n_0_72), .Q(\r_values[0] [15]), 
      .QN());
   DFF_X1 \r_values_reg[0][14]  (.D(n_0_51), .CK(n_0_72), .Q(\r_values[0] [14]), 
      .QN());
   DFF_X1 \r_values_reg[0][13]  (.D(n_0_52), .CK(n_0_72), .Q(\r_values[0] [13]), 
      .QN());
   DFF_X1 \r_values_reg[0][12]  (.D(n_0_53), .CK(n_0_72), .Q(\r_values[0] [12]), 
      .QN());
   DFF_X1 \r_values_reg[0][11]  (.D(n_0_54), .CK(n_0_72), .Q(\r_values[0] [11]), 
      .QN());
   DFF_X1 \r_values_reg[0][10]  (.D(n_0_55), .CK(n_0_72), .Q(\r_values[0] [10]), 
      .QN());
   DFF_X1 \r_values_reg[0][9]  (.D(n_0_56), .CK(n_0_72), .Q(\r_values[0] [9]), 
      .QN());
   DFF_X1 \r_values_reg[0][8]  (.D(n_0_57), .CK(n_0_72), .Q(\r_values[0] [8]), 
      .QN());
   DFF_X1 \r_values_reg[0][7]  (.D(n_0_58), .CK(n_0_72), .Q(\r_values[0] [7]), 
      .QN());
   DFF_X1 \r_values_reg[0][6]  (.D(n_0_59), .CK(n_0_72), .Q(\r_values[0] [6]), 
      .QN());
   DFF_X1 \r_values_reg[0][5]  (.D(n_0_60), .CK(n_0_72), .Q(\r_values[0] [5]), 
      .QN());
   DFF_X1 \r_values_reg[0][4]  (.D(n_0_61), .CK(n_0_72), .Q(\r_values[0] [4]), 
      .QN());
   DFF_X1 \r_values_reg[0][3]  (.D(n_0_62), .CK(n_0_72), .Q(\r_values[0] [3]), 
      .QN());
   DFF_X1 \r_values_reg[0][2]  (.D(n_0_63), .CK(n_0_72), .Q(\r_values[0] [2]), 
      .QN());
   DFF_X1 \r_values_reg[0][1]  (.D(n_0_64), .CK(n_0_72), .Q(\r_values[0] [1]), 
      .QN());
   DFF_X1 \r_values_reg[0][0]  (.D(n_0_65), .CK(n_0_72), .Q(\r_values[0] [0]), 
      .QN());
   DFF_X1 \r_values_reg[1][15]  (.D(n_0_66), .CK(n_0_72), .Q(\r_values[1] [15]), 
      .QN());
   DFF_X1 \r_values_reg[1][14]  (.D(n_0_67), .CK(n_0_72), .Q(\r_values[1] [14]), 
      .QN());
   DFF_X1 \r_values_reg[1][13]  (.D(n_0_68), .CK(n_0_72), .Q(\r_values[1] [13]), 
      .QN());
   DFF_X1 \r_values_reg[1][12]  (.D(n_0_69), .CK(n_0_72), .Q(\r_values[1] [12]), 
      .QN());
   DFF_X1 \r_values_reg[1][11]  (.D(n_0_70), .CK(n_0_72), .Q(\r_values[1] [11]), 
      .QN());
   DFF_X1 \r_values_reg[1][10]  (.D(n_0_71), .CK(n_0_72), .Q(\r_values[1] [10]), 
      .QN());
   DFF_X1 \r_values_reg[1][9]  (.D(n_0_73), .CK(n_0_72), .Q(\r_values[1] [9]), 
      .QN());
   DFF_X1 \r_values_reg[1][8]  (.D(n_0_74), .CK(n_0_72), .Q(\r_values[1] [8]), 
      .QN());
   DFF_X1 \r_values_reg[1][7]  (.D(n_0_75), .CK(n_0_72), .Q(\r_values[1] [7]), 
      .QN());
   DFF_X1 \r_values_reg[1][6]  (.D(n_0_76), .CK(n_0_72), .Q(\r_values[1] [6]), 
      .QN());
   DFF_X1 \r_values_reg[1][5]  (.D(n_0_77), .CK(n_0_72), .Q(\r_values[1] [5]), 
      .QN());
   DFF_X1 \r_values_reg[1][4]  (.D(n_0_78), .CK(n_0_72), .Q(\r_values[1] [4]), 
      .QN());
   DFF_X1 \r_values_reg[1][3]  (.D(n_0_79), .CK(n_0_72), .Q(\r_values[1] [3]), 
      .QN());
   DFF_X1 \r_values_reg[1][2]  (.D(n_0_80), .CK(n_0_72), .Q(\r_values[1] [2]), 
      .QN());
   DFF_X1 \r_values_reg[1][1]  (.D(n_0_49), .CK(n_0_72), .Q(\r_values[1] [1]), 
      .QN());
   DFF_X1 \r_values_reg[1][0]  (.D(n_0_48), .CK(n_0_72), .Q(\r_values[1] [0]), 
      .QN());
   DFF_X1 \r_weights_reg[0][15]  (.D(n_0_47), .CK(n_0_72), .Q(\r_weights[0] [15]), 
      .QN());
   DFF_X1 \r_weights_reg[0][14]  (.D(n_0_46), .CK(n_0_72), .Q(\r_weights[0] [14]), 
      .QN());
   DFF_X1 \r_weights_reg[0][13]  (.D(n_0_45), .CK(n_0_72), .Q(\r_weights[0] [13]), 
      .QN());
   DFF_X1 \r_weights_reg[0][12]  (.D(n_0_44), .CK(n_0_72), .Q(\r_weights[0] [12]), 
      .QN());
   DFF_X1 \r_weights_reg[0][11]  (.D(n_0_43), .CK(n_0_72), .Q(\r_weights[0] [11]), 
      .QN());
   DFF_X1 \r_weights_reg[0][10]  (.D(n_0_42), .CK(n_0_72), .Q(\r_weights[0] [10]), 
      .QN());
   DFF_X1 \r_weights_reg[0][9]  (.D(n_0_41), .CK(n_0_72), .Q(\r_weights[0] [9]), 
      .QN());
   DFF_X1 \r_weights_reg[0][8]  (.D(n_0_40), .CK(n_0_72), .Q(\r_weights[0] [8]), 
      .QN());
   DFF_X1 \r_weights_reg[0][7]  (.D(n_0_39), .CK(n_0_72), .Q(\r_weights[0] [7]), 
      .QN());
   DFF_X1 \r_weights_reg[0][6]  (.D(n_0_38), .CK(n_0_72), .Q(\r_weights[0] [6]), 
      .QN());
   DFF_X1 \r_weights_reg[0][5]  (.D(n_0_37), .CK(n_0_72), .Q(\r_weights[0] [5]), 
      .QN());
   DFF_X1 \r_weights_reg[0][4]  (.D(n_0_36), .CK(n_0_72), .Q(\r_weights[0] [4]), 
      .QN());
   DFF_X1 \r_weights_reg[0][3]  (.D(n_0_35), .CK(n_0_72), .Q(\r_weights[0] [3]), 
      .QN());
   DFF_X1 \r_weights_reg[0][2]  (.D(n_0_34), .CK(n_0_72), .Q(\r_weights[0] [2]), 
      .QN());
   DFF_X1 \r_weights_reg[0][1]  (.D(n_0_33), .CK(n_0_72), .Q(\r_weights[0] [1]), 
      .QN());
   DFF_X1 \r_weights_reg[0][0]  (.D(n_0_32), .CK(n_0_72), .Q(\r_weights[0] [0]), 
      .QN());
   DFF_X1 \r_weights_reg[1][15]  (.D(n_0_31), .CK(n_0_72), .Q(\r_weights[1] [15]), 
      .QN());
   DFF_X1 \r_weights_reg[1][14]  (.D(n_0_30), .CK(n_0_72), .Q(\r_weights[1] [14]), 
      .QN());
   DFF_X1 \r_weights_reg[1][13]  (.D(n_0_29), .CK(n_0_72), .Q(\r_weights[1] [13]), 
      .QN());
   DFF_X1 \r_weights_reg[1][12]  (.D(n_0_28), .CK(n_0_72), .Q(\r_weights[1] [12]), 
      .QN());
   DFF_X1 \r_weights_reg[1][11]  (.D(n_0_27), .CK(n_0_72), .Q(\r_weights[1] [11]), 
      .QN());
   DFF_X1 \r_weights_reg[1][10]  (.D(n_0_26), .CK(n_0_72), .Q(\r_weights[1] [10]), 
      .QN());
   DFF_X1 \r_weights_reg[1][9]  (.D(n_0_25), .CK(n_0_72), .Q(\r_weights[1] [9]), 
      .QN());
   DFF_X1 \r_weights_reg[1][8]  (.D(n_0_24), .CK(n_0_72), .Q(\r_weights[1] [8]), 
      .QN());
   DFF_X1 \r_weights_reg[1][7]  (.D(n_0_23), .CK(n_0_72), .Q(\r_weights[1] [7]), 
      .QN());
   DFF_X1 \r_weights_reg[1][6]  (.D(n_0_22), .CK(n_0_72), .Q(\r_weights[1] [6]), 
      .QN());
   DFF_X1 \r_weights_reg[1][5]  (.D(n_0_21), .CK(n_0_72), .Q(\r_weights[1] [5]), 
      .QN());
   DFF_X1 \r_weights_reg[1][4]  (.D(n_0_20), .CK(n_0_72), .Q(\r_weights[1] [4]), 
      .QN());
   DFF_X1 \r_weights_reg[1][3]  (.D(n_0_19), .CK(n_0_72), .Q(\r_weights[1] [3]), 
      .QN());
   DFF_X1 \r_weights_reg[1][2]  (.D(n_0_18), .CK(n_0_72), .Q(\r_weights[1] [2]), 
      .QN());
   DFF_X1 \r_weights_reg[1][1]  (.D(n_0_17), .CK(n_0_72), .Q(\r_weights[1] [1]), 
      .QN());
   DFF_X1 \r_weights_reg[1][0]  (.D(n_0_16), .CK(n_0_72), .Q(\r_weights[1] [0]), 
      .QN());
   DFF_X1 \r_bias_reg[15]  (.D(n_0_15), .CK(n_0_72), .Q(r_bias[15]), .QN());
   DFF_X1 \r_bias_reg[14]  (.D(n_0_14), .CK(n_0_72), .Q(r_bias[14]), .QN());
   DFF_X1 \r_bias_reg[13]  (.D(n_0_13), .CK(n_0_72), .Q(r_bias[13]), .QN());
   DFF_X1 \r_bias_reg[12]  (.D(n_0_12), .CK(n_0_72), .Q(r_bias[12]), .QN());
   DFF_X1 \r_bias_reg[11]  (.D(n_0_11), .CK(n_0_72), .Q(r_bias[11]), .QN());
   DFF_X1 \r_bias_reg[10]  (.D(n_0_10), .CK(n_0_72), .Q(r_bias[10]), .QN());
   DFF_X1 \r_bias_reg[9]  (.D(n_0_9), .CK(n_0_72), .Q(r_bias[9]), .QN());
   DFF_X1 \r_bias_reg[8]  (.D(n_0_8), .CK(n_0_72), .Q(r_bias[8]), .QN());
   DFF_X1 \r_bias_reg[7]  (.D(n_0_7), .CK(n_0_72), .Q(r_bias[7]), .QN());
   DFF_X1 \r_bias_reg[6]  (.D(n_0_6), .CK(n_0_72), .Q(r_bias[6]), .QN());
   DFF_X1 \r_bias_reg[5]  (.D(n_0_5), .CK(n_0_72), .Q(r_bias[5]), .QN());
   DFF_X1 \r_bias_reg[4]  (.D(n_0_4), .CK(n_0_72), .Q(r_bias[4]), .QN());
   DFF_X1 \r_bias_reg[3]  (.D(n_0_3), .CK(n_0_72), .Q(r_bias[3]), .QN());
   DFF_X1 \r_bias_reg[2]  (.D(n_0_2), .CK(n_0_72), .Q(r_bias[2]), .QN());
   DFF_X1 \r_bias_reg[1]  (.D(n_0_1), .CK(n_0_72), .Q(r_bias[1]), .QN());
   DFF_X1 \r_bias_reg[0]  (.D(n_0_0), .CK(n_0_72), .Q(r_bias[0]), .QN());
   INV_X1 i_0_1_0 (.A(n_0_1_0), .ZN(n_0_0));
   AOI22_X1 i_0_1_1 (.A1(i_single[0]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[0]), .ZN(n_0_1_0));
   INV_X1 i_0_1_2 (.A(n_0_1_1), .ZN(n_0_1));
   AOI22_X1 i_0_1_3 (.A1(i_single[1]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[1]), .ZN(n_0_1_1));
   INV_X1 i_0_1_4 (.A(n_0_1_2), .ZN(n_0_2));
   AOI22_X1 i_0_1_5 (.A1(i_single[2]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[2]), .ZN(n_0_1_2));
   INV_X1 i_0_1_6 (.A(n_0_1_3), .ZN(n_0_3));
   AOI22_X1 i_0_1_7 (.A1(i_single[3]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[3]), .ZN(n_0_1_3));
   INV_X1 i_0_1_8 (.A(n_0_1_4), .ZN(n_0_4));
   AOI22_X1 i_0_1_9 (.A1(i_single[4]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[4]), .ZN(n_0_1_4));
   INV_X1 i_0_1_10 (.A(n_0_1_5), .ZN(n_0_5));
   AOI22_X1 i_0_1_11 (.A1(i_single[5]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[5]), .ZN(n_0_1_5));
   INV_X1 i_0_1_12 (.A(n_0_1_6), .ZN(n_0_6));
   AOI22_X1 i_0_1_13 (.A1(i_single[6]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[6]), .ZN(n_0_1_6));
   INV_X1 i_0_1_14 (.A(n_0_1_7), .ZN(n_0_7));
   AOI22_X1 i_0_1_15 (.A1(i_single[7]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[7]), .ZN(n_0_1_7));
   INV_X1 i_0_1_16 (.A(n_0_1_8), .ZN(n_0_8));
   AOI22_X1 i_0_1_17 (.A1(i_single[8]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[8]), .ZN(n_0_1_8));
   INV_X1 i_0_1_18 (.A(n_0_1_9), .ZN(n_0_9));
   AOI22_X1 i_0_1_19 (.A1(i_single[9]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[9]), .ZN(n_0_1_9));
   INV_X1 i_0_1_20 (.A(n_0_1_10), .ZN(n_0_10));
   AOI22_X1 i_0_1_21 (.A1(i_single[10]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[10]), .ZN(n_0_1_10));
   INV_X1 i_0_1_22 (.A(n_0_1_11), .ZN(n_0_11));
   AOI22_X1 i_0_1_23 (.A1(i_single[11]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[11]), .ZN(n_0_1_11));
   INV_X1 i_0_1_24 (.A(n_0_1_12), .ZN(n_0_12));
   AOI22_X1 i_0_1_25 (.A1(i_single[12]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[12]), .ZN(n_0_1_12));
   INV_X1 i_0_1_26 (.A(n_0_1_13), .ZN(n_0_13));
   AOI22_X1 i_0_1_27 (.A1(i_single[13]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[13]), .ZN(n_0_1_13));
   INV_X1 i_0_1_28 (.A(n_0_1_14), .ZN(n_0_14));
   AOI22_X1 i_0_1_29 (.A1(i_single[14]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[14]), .ZN(n_0_1_14));
   INV_X1 i_0_1_30 (.A(n_0_1_15), .ZN(n_0_15));
   AOI22_X1 i_0_1_31 (.A1(i_single[15]), .A2(n_0_1_49), .B1(n_0_1_48), .B2(
      r_bias[15]), .ZN(n_0_1_15));
   INV_X1 i_0_1_32 (.A(n_0_1_16), .ZN(n_0_16));
   AOI22_X1 i_0_1_33 (.A1(\i_values[1] [0]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [0]), .ZN(n_0_1_16));
   INV_X1 i_0_1_34 (.A(n_0_1_17), .ZN(n_0_17));
   AOI22_X1 i_0_1_35 (.A1(\i_values[1] [1]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [1]), .ZN(n_0_1_17));
   INV_X1 i_0_1_36 (.A(n_0_1_18), .ZN(n_0_18));
   AOI22_X1 i_0_1_37 (.A1(\i_values[1] [2]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [2]), .ZN(n_0_1_18));
   INV_X1 i_0_1_38 (.A(n_0_1_19), .ZN(n_0_19));
   AOI22_X1 i_0_1_39 (.A1(\i_values[1] [3]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [3]), .ZN(n_0_1_19));
   INV_X1 i_0_1_40 (.A(n_0_1_20), .ZN(n_0_20));
   AOI22_X1 i_0_1_41 (.A1(\i_values[1] [4]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [4]), .ZN(n_0_1_20));
   INV_X1 i_0_1_42 (.A(n_0_1_21), .ZN(n_0_21));
   AOI22_X1 i_0_1_43 (.A1(\i_values[1] [5]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [5]), .ZN(n_0_1_21));
   INV_X1 i_0_1_44 (.A(n_0_1_22), .ZN(n_0_22));
   AOI22_X1 i_0_1_45 (.A1(\i_values[1] [6]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [6]), .ZN(n_0_1_22));
   INV_X1 i_0_1_46 (.A(n_0_1_23), .ZN(n_0_23));
   AOI22_X1 i_0_1_47 (.A1(\i_values[1] [7]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [7]), .ZN(n_0_1_23));
   INV_X1 i_0_1_48 (.A(n_0_1_24), .ZN(n_0_24));
   AOI22_X1 i_0_1_49 (.A1(\i_values[1] [8]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [8]), .ZN(n_0_1_24));
   INV_X1 i_0_1_50 (.A(n_0_1_25), .ZN(n_0_25));
   AOI22_X1 i_0_1_51 (.A1(\i_values[1] [9]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [9]), .ZN(n_0_1_25));
   INV_X1 i_0_1_52 (.A(n_0_1_26), .ZN(n_0_26));
   AOI22_X1 i_0_1_53 (.A1(\i_values[1] [10]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [10]), .ZN(n_0_1_26));
   INV_X1 i_0_1_54 (.A(n_0_1_27), .ZN(n_0_27));
   AOI22_X1 i_0_1_55 (.A1(\i_values[1] [11]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [11]), .ZN(n_0_1_27));
   INV_X1 i_0_1_56 (.A(n_0_1_28), .ZN(n_0_28));
   AOI22_X1 i_0_1_57 (.A1(\i_values[1] [12]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [12]), .ZN(n_0_1_28));
   INV_X1 i_0_1_58 (.A(n_0_1_29), .ZN(n_0_29));
   AOI22_X1 i_0_1_59 (.A1(\i_values[1] [13]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [13]), .ZN(n_0_1_29));
   INV_X1 i_0_1_60 (.A(n_0_1_30), .ZN(n_0_30));
   AOI22_X1 i_0_1_61 (.A1(\i_values[1] [14]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [14]), .ZN(n_0_1_30));
   INV_X1 i_0_1_62 (.A(n_0_1_31), .ZN(n_0_31));
   AOI22_X1 i_0_1_63 (.A1(\i_values[1] [15]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[1] [15]), .ZN(n_0_1_31));
   INV_X1 i_0_1_64 (.A(n_0_1_32), .ZN(n_0_32));
   AOI22_X1 i_0_1_65 (.A1(\i_values[0] [0]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [0]), .ZN(n_0_1_32));
   INV_X1 i_0_1_66 (.A(n_0_1_33), .ZN(n_0_33));
   AOI22_X1 i_0_1_67 (.A1(\i_values[0] [1]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [1]), .ZN(n_0_1_33));
   INV_X1 i_0_1_68 (.A(n_0_1_34), .ZN(n_0_34));
   AOI22_X1 i_0_1_69 (.A1(\i_values[0] [2]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [2]), .ZN(n_0_1_34));
   INV_X1 i_0_1_70 (.A(n_0_1_35), .ZN(n_0_35));
   AOI22_X1 i_0_1_71 (.A1(\i_values[0] [3]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [3]), .ZN(n_0_1_35));
   INV_X1 i_0_1_72 (.A(n_0_1_36), .ZN(n_0_36));
   AOI22_X1 i_0_1_73 (.A1(\i_values[0] [4]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [4]), .ZN(n_0_1_36));
   INV_X1 i_0_1_74 (.A(n_0_1_37), .ZN(n_0_37));
   AOI22_X1 i_0_1_75 (.A1(\i_values[0] [5]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [5]), .ZN(n_0_1_37));
   INV_X1 i_0_1_76 (.A(n_0_1_38), .ZN(n_0_38));
   AOI22_X1 i_0_1_77 (.A1(\i_values[0] [6]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [6]), .ZN(n_0_1_38));
   INV_X1 i_0_1_78 (.A(n_0_1_39), .ZN(n_0_39));
   AOI22_X1 i_0_1_79 (.A1(\i_values[0] [7]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [7]), .ZN(n_0_1_39));
   INV_X1 i_0_1_80 (.A(n_0_1_40), .ZN(n_0_40));
   AOI22_X1 i_0_1_81 (.A1(\i_values[0] [8]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [8]), .ZN(n_0_1_40));
   INV_X1 i_0_1_82 (.A(n_0_1_41), .ZN(n_0_41));
   AOI22_X1 i_0_1_83 (.A1(\i_values[0] [9]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [9]), .ZN(n_0_1_41));
   INV_X1 i_0_1_84 (.A(n_0_1_42), .ZN(n_0_42));
   AOI22_X1 i_0_1_85 (.A1(\i_values[0] [10]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [10]), .ZN(n_0_1_42));
   INV_X1 i_0_1_86 (.A(n_0_1_43), .ZN(n_0_43));
   AOI22_X1 i_0_1_87 (.A1(\i_values[0] [11]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [11]), .ZN(n_0_1_43));
   INV_X1 i_0_1_88 (.A(n_0_1_44), .ZN(n_0_44));
   AOI22_X1 i_0_1_89 (.A1(\i_values[0] [12]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [12]), .ZN(n_0_1_44));
   INV_X1 i_0_1_90 (.A(n_0_1_45), .ZN(n_0_45));
   AOI22_X1 i_0_1_91 (.A1(\i_values[0] [13]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [13]), .ZN(n_0_1_45));
   INV_X1 i_0_1_92 (.A(n_0_1_46), .ZN(n_0_46));
   AOI22_X1 i_0_1_93 (.A1(\i_values[0] [14]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [14]), .ZN(n_0_1_46));
   INV_X1 i_0_1_94 (.A(n_0_1_47), .ZN(n_0_47));
   AOI22_X1 i_0_1_95 (.A1(\i_values[0] [15]), .A2(n_0_1_49), .B1(n_0_1_48), 
      .B2(\r_weights[0] [15]), .ZN(n_0_1_47));
   AOI21_X1 i_0_1_96 (.A(clear), .B1(n_0_1_52), .B2(load_enable[0]), .ZN(
      n_0_1_48));
   NOR3_X1 i_0_1_97 (.A1(n_0_1_51), .A2(load_enable[1]), .A3(clear), .ZN(
      n_0_1_49));
   MUX2_X1 i_0_1_98 (.A(\i_values[1] [0]), .B(\r_values[1] [0]), .S(n_0_1_50), 
      .Z(n_0_48));
   MUX2_X1 i_0_1_99 (.A(\i_values[1] [1]), .B(\r_values[1] [1]), .S(n_0_1_50), 
      .Z(n_0_49));
   MUX2_X1 i_0_1_100 (.A(\i_values[1] [2]), .B(\r_values[1] [2]), .S(n_0_1_50), 
      .Z(n_0_80));
   MUX2_X1 i_0_1_101 (.A(\i_values[1] [3]), .B(\r_values[1] [3]), .S(n_0_1_50), 
      .Z(n_0_79));
   MUX2_X1 i_0_1_102 (.A(\i_values[1] [4]), .B(\r_values[1] [4]), .S(n_0_1_50), 
      .Z(n_0_78));
   MUX2_X1 i_0_1_103 (.A(\i_values[1] [5]), .B(\r_values[1] [5]), .S(n_0_1_50), 
      .Z(n_0_77));
   MUX2_X1 i_0_1_104 (.A(\i_values[1] [6]), .B(\r_values[1] [6]), .S(n_0_1_50), 
      .Z(n_0_76));
   MUX2_X1 i_0_1_105 (.A(\i_values[1] [7]), .B(\r_values[1] [7]), .S(n_0_1_50), 
      .Z(n_0_75));
   MUX2_X1 i_0_1_106 (.A(\i_values[1] [8]), .B(\r_values[1] [8]), .S(n_0_1_50), 
      .Z(n_0_74));
   MUX2_X1 i_0_1_107 (.A(\i_values[1] [9]), .B(\r_values[1] [9]), .S(n_0_1_50), 
      .Z(n_0_73));
   MUX2_X1 i_0_1_108 (.A(\i_values[1] [10]), .B(\r_values[1] [10]), .S(n_0_1_50), 
      .Z(n_0_71));
   MUX2_X1 i_0_1_109 (.A(\i_values[1] [11]), .B(\r_values[1] [11]), .S(n_0_1_50), 
      .Z(n_0_70));
   MUX2_X1 i_0_1_110 (.A(\i_values[1] [12]), .B(\r_values[1] [12]), .S(n_0_1_50), 
      .Z(n_0_69));
   MUX2_X1 i_0_1_111 (.A(\i_values[1] [13]), .B(\r_values[1] [13]), .S(n_0_1_50), 
      .Z(n_0_68));
   MUX2_X1 i_0_1_112 (.A(\i_values[1] [14]), .B(\r_values[1] [14]), .S(n_0_1_50), 
      .Z(n_0_67));
   MUX2_X1 i_0_1_113 (.A(\i_values[1] [15]), .B(\r_values[1] [15]), .S(n_0_1_50), 
      .Z(n_0_66));
   MUX2_X1 i_0_1_114 (.A(\i_values[0] [0]), .B(\r_values[0] [0]), .S(n_0_1_50), 
      .Z(n_0_65));
   MUX2_X1 i_0_1_115 (.A(\i_values[0] [1]), .B(\r_values[0] [1]), .S(n_0_1_50), 
      .Z(n_0_64));
   MUX2_X1 i_0_1_116 (.A(\i_values[0] [2]), .B(\r_values[0] [2]), .S(n_0_1_50), 
      .Z(n_0_63));
   MUX2_X1 i_0_1_117 (.A(\i_values[0] [3]), .B(\r_values[0] [3]), .S(n_0_1_50), 
      .Z(n_0_62));
   MUX2_X1 i_0_1_118 (.A(\i_values[0] [4]), .B(\r_values[0] [4]), .S(n_0_1_50), 
      .Z(n_0_61));
   MUX2_X1 i_0_1_119 (.A(\i_values[0] [5]), .B(\r_values[0] [5]), .S(n_0_1_50), 
      .Z(n_0_60));
   MUX2_X1 i_0_1_120 (.A(\i_values[0] [6]), .B(\r_values[0] [6]), .S(n_0_1_50), 
      .Z(n_0_59));
   MUX2_X1 i_0_1_121 (.A(\i_values[0] [7]), .B(\r_values[0] [7]), .S(n_0_1_50), 
      .Z(n_0_58));
   MUX2_X1 i_0_1_122 (.A(\i_values[0] [8]), .B(\r_values[0] [8]), .S(n_0_1_50), 
      .Z(n_0_57));
   MUX2_X1 i_0_1_123 (.A(\i_values[0] [9]), .B(\r_values[0] [9]), .S(n_0_1_50), 
      .Z(n_0_56));
   MUX2_X1 i_0_1_124 (.A(\i_values[0] [10]), .B(\r_values[0] [10]), .S(n_0_1_50), 
      .Z(n_0_55));
   MUX2_X1 i_0_1_125 (.A(\i_values[0] [11]), .B(\r_values[0] [11]), .S(n_0_1_50), 
      .Z(n_0_54));
   MUX2_X1 i_0_1_126 (.A(\i_values[0] [12]), .B(\r_values[0] [12]), .S(n_0_1_50), 
      .Z(n_0_53));
   MUX2_X1 i_0_1_127 (.A(\i_values[0] [13]), .B(\r_values[0] [13]), .S(n_0_1_50), 
      .Z(n_0_52));
   MUX2_X1 i_0_1_128 (.A(\i_values[0] [14]), .B(\r_values[0] [14]), .S(n_0_1_50), 
      .Z(n_0_51));
   MUX2_X1 i_0_1_129 (.A(\i_values[0] [15]), .B(\r_values[0] [15]), .S(n_0_1_50), 
      .Z(n_0_50));
   OR3_X1 i_0_1_130 (.A1(clear), .A2(load_enable[1]), .A3(load_enable[0]), 
      .ZN(n_0_1_50));
   INV_X1 i_0_1_131 (.A(load_enable[0]), .ZN(n_0_1_51));
   INV_X1 i_0_1_132 (.A(load_enable[1]), .ZN(n_0_1_52));
   INV_X1 i_0_1_133 (.A(clk), .ZN(n_0_72));
endmodule
