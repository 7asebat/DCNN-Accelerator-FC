
// 	Thu May  6 06:06:25 2021
//	vlsi
//	localhost.localdomain

module Neuron_Layer (clk, load_en, load_value, load_address, reset, \values[0] , 
    \values[1] , \values[2] , \values[3] , \values[4] , \values[5] , \values[6] , 
    \values[7] , \values[8] , \values[9] , \values[10] , \values[11] , \values[12] , 
    \values[13] , \values[14] , \values[15] , \values[16] , \values[17] , \values[18] , 
    \values[19] , \values[20] , \values[21] , \values[22] , \values[23] , \values[24] , 
    \values[25] , \values[26] , \values[27] , \values[28] , \values[29] , \values[30] , 
    \values[31] , \values[32] , \values[33] , \values[34] , \values[35] , \values[36] , 
    \values[37] , \values[38] , \values[39] , \values[40] , \values[41] , \values[42] , 
    \values[43] , \values[44] , \values[45] , \values[46] , \values[47] , \values[48] , 
    \values[49] , \values[50] , \values[51] , \values[52] , \values[53] , \values[54] , 
    \values[55] , \values[56] , \values[57] , \values[58] , \values[59] , \values[60] , 
    \values[61] , \values[62] , \values[63] , \values[64] , \values[65] , \values[66] , 
    \values[67] , \values[68] , \values[69] , \values[70] , \values[71] , \values[72] , 
    \values[73] , \values[74] , \values[75] , \values[76] , \values[77] , \values[78] , 
    \values[79] , \values[80] , \values[81] , \values[82] , \values[83] , \values[84] , 
    \values[85] , \values[86] , \values[87] , \values[88] , \values[89] , \values[90] , 
    \values[91] , \values[92] , \values[93] , \values[94] , \values[95] , \values[96] , 
    \values[97] , \values[98] , \values[99] , \values[100] , \values[101] , \values[102] , 
    \values[103] , \values[104] , \values[105] , \values[106] , \values[107] , \values[108] , 
    \values[109] , \values[110] , \values[111] , \values[112] , \values[113] , \values[114] , 
    \values[115] , \values[116] , \values[117] , \values[118] , \values[119] );

output [15:0] \values[0] ;
output [15:0] \values[100] ;
output [15:0] \values[101] ;
output [15:0] \values[102] ;
output [15:0] \values[103] ;
output [15:0] \values[104] ;
output [15:0] \values[105] ;
output [15:0] \values[106] ;
output [15:0] \values[107] ;
output [15:0] \values[108] ;
output [15:0] \values[109] ;
output [15:0] \values[10] ;
output [15:0] \values[110] ;
output [15:0] \values[111] ;
output [15:0] \values[112] ;
output [15:0] \values[113] ;
output [15:0] \values[114] ;
output [15:0] \values[115] ;
output [15:0] \values[116] ;
output [15:0] \values[117] ;
output [15:0] \values[118] ;
output [15:0] \values[119] ;
output [15:0] \values[11] ;
output [15:0] \values[12] ;
output [15:0] \values[13] ;
output [15:0] \values[14] ;
output [15:0] \values[15] ;
output [15:0] \values[16] ;
output [15:0] \values[17] ;
output [15:0] \values[18] ;
output [15:0] \values[19] ;
output [15:0] \values[1] ;
output [15:0] \values[20] ;
output [15:0] \values[21] ;
output [15:0] \values[22] ;
output [15:0] \values[23] ;
output [15:0] \values[24] ;
output [15:0] \values[25] ;
output [15:0] \values[26] ;
output [15:0] \values[27] ;
output [15:0] \values[28] ;
output [15:0] \values[29] ;
output [15:0] \values[2] ;
output [15:0] \values[30] ;
output [15:0] \values[31] ;
output [15:0] \values[32] ;
output [15:0] \values[33] ;
output [15:0] \values[34] ;
output [15:0] \values[35] ;
output [15:0] \values[36] ;
output [15:0] \values[37] ;
output [15:0] \values[38] ;
output [15:0] \values[39] ;
output [15:0] \values[3] ;
output [15:0] \values[40] ;
output [15:0] \values[41] ;
output [15:0] \values[42] ;
output [15:0] \values[43] ;
output [15:0] \values[44] ;
output [15:0] \values[45] ;
output [15:0] \values[46] ;
output [15:0] \values[47] ;
output [15:0] \values[48] ;
output [15:0] \values[49] ;
output [15:0] \values[4] ;
output [15:0] \values[50] ;
output [15:0] \values[51] ;
output [15:0] \values[52] ;
output [15:0] \values[53] ;
output [15:0] \values[54] ;
output [15:0] \values[55] ;
output [15:0] \values[56] ;
output [15:0] \values[57] ;
output [15:0] \values[58] ;
output [15:0] \values[59] ;
output [15:0] \values[5] ;
output [15:0] \values[60] ;
output [15:0] \values[61] ;
output [15:0] \values[62] ;
output [15:0] \values[63] ;
output [15:0] \values[64] ;
output [15:0] \values[65] ;
output [15:0] \values[66] ;
output [15:0] \values[67] ;
output [15:0] \values[68] ;
output [15:0] \values[69] ;
output [15:0] \values[6] ;
output [15:0] \values[70] ;
output [15:0] \values[71] ;
output [15:0] \values[72] ;
output [15:0] \values[73] ;
output [15:0] \values[74] ;
output [15:0] \values[75] ;
output [15:0] \values[76] ;
output [15:0] \values[77] ;
output [15:0] \values[78] ;
output [15:0] \values[79] ;
output [15:0] \values[7] ;
output [15:0] \values[80] ;
output [15:0] \values[81] ;
output [15:0] \values[82] ;
output [15:0] \values[83] ;
output [15:0] \values[84] ;
output [15:0] \values[85] ;
output [15:0] \values[86] ;
output [15:0] \values[87] ;
output [15:0] \values[88] ;
output [15:0] \values[89] ;
output [15:0] \values[8] ;
output [15:0] \values[90] ;
output [15:0] \values[91] ;
output [15:0] \values[92] ;
output [15:0] \values[93] ;
output [15:0] \values[94] ;
output [15:0] \values[95] ;
output [15:0] \values[96] ;
output [15:0] \values[97] ;
output [15:0] \values[98] ;
output [15:0] \values[99] ;
output [15:0] \values[9] ;
input clk;
input [15:0] load_address;
input load_en;
input [15:0] load_value;
input reset;
wire n_121_0;
wire n_121_1;
wire n_121_2;
wire n_121_3;
wire n_121_4;
wire n_121_5;
wire n_121_6;
wire n_121_7;
wire n_121_8;
wire n_121_9;
wire n_121_10;
wire n_121_11;
wire n_121_12;
wire n_121_13;
wire n_121_14;
wire n_121_15;
wire n_121_16;
wire n_121_17;
wire n_121_18;
wire n_121_19;
wire n_121_20;
wire n_121_21;
wire n_121_22;
wire n_121_23;
wire n_121_24;
wire n_121_25;
wire n_121_26;
wire n_121_27;
wire n_121_28;
wire n_121_29;
wire n_121_30;
wire n_121_31;
wire n_121_32;
wire n_121_33;
wire n_121_34;
wire n_121_35;
wire n_121_36;
wire n_121_37;
wire n_121_38;
wire n_121_39;
wire n_121_40;
wire n_121_41;
wire n_121_42;
wire n_121_43;
wire n_121_44;
wire n_121_45;
wire n_121_46;
wire n_121_47;
wire n_121_48;
wire n_121_49;
wire n_121_50;
wire n_121_51;
wire n_121_52;
wire n_121_53;
wire n_121_54;
wire n_121_55;
wire n_121_56;
wire n_121_57;
wire n_121_58;
wire n_121_59;
wire n_121_60;
wire n_121_61;
wire n_121_62;
wire n_121_63;
wire n_121_64;
wire n_121_65;
wire n_121_66;
wire n_121_67;
wire n_121_68;
wire n_121_69;
wire n_121_70;
wire n_121_71;
wire n_121_72;
wire n_121_73;
wire n_121_74;
wire n_121_75;
wire n_121_76;
wire n_121_77;
wire n_121_78;
wire n_121_79;
wire n_121_80;
wire n_121_81;
wire n_121_82;
wire n_121_83;
wire n_121_84;
wire n_121_85;
wire n_121_86;
wire n_121_87;
wire n_121_88;
wire n_121_89;
wire n_121_90;
wire n_121_91;
wire n_121_92;
wire n_121_93;
wire n_122_0;
wire n_122_1;
wire n_122_2;
wire n_122_3;
wire n_122_4;
wire n_122_5;
wire n_122_6;
wire n_122_7;
wire n_122_8;
wire n_122_9;
wire n_122_10;
wire n_122_11;
wire n_122_12;
wire n_122_13;
wire n_122_14;
wire n_122_15;
wire n_122_16;
wire n_122_17;
wire n_122_18;
wire n_122_19;
wire n_122_20;
wire n_122_21;
wire n_122_22;
wire n_122_23;
wire n_122_24;
wire n_122_25;
wire n_0_0_0;
wire \values[15] ;
wire \values[14] ;
wire \values[13] ;
wire \values[12] ;
wire \values[11] ;
wire \values[10] ;
wire \values[9] ;
wire \values[8] ;
wire \values[7] ;
wire \values[6] ;
wire \values[5] ;
wire \values[4] ;
wire \values[3] ;
wire \values[2] ;
wire \values[1] ;
wire \values[0] ;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_96;
wire n_95;
wire n_94;
wire n_93;
wire n_92;
wire n_91;
wire n_90;
wire n_89;
wire n_88;
wire n_87;
wire n_86;
wire n_85;
wire n_84;
wire n_83;
wire n_82;
wire n_81;
wire n_80;
wire n_79;
wire n_78;
wire n_77;
wire n_76;
wire n_75;
wire n_74;
wire n_73;
wire n_72;
wire n_71;
wire n_70;
wire n_69;
wire n_68;
wire n_67;
wire n_66;
wire n_65;
wire n_64;
wire n_63;
wire n_62;
wire n_61;
wire n_60;
wire n_59;
wire n_58;
wire n_57;
wire n_56;
wire n_55;
wire n_54;
wire n_53;
wire n_52;
wire n_51;
wire n_50;
wire n_49;
wire n_48;
wire n_47;
wire n_46;
wire n_45;
wire n_44;
wire n_43;
wire n_42;
wire n_41;
wire n_40;
wire n_39;
wire n_38;
wire n_37;
wire n_36;
wire n_35;
wire n_34;
wire n_33;
wire n_32;
wire n_31;
wire n_30;
wire n_29;
wire n_28;
wire n_27;
wire n_26;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_2;
wire n_1;
wire n_0;
wire sps__n1;
wire sps__n4;
wire sps__n5;
wire sps__n10;
wire sps__n11;
wire sps__n12;
wire spc__n157;
wire sps__n14;
wire sps__n25;
wire spc__n158;
wire sps__n27;
wire sps__n28;
wire sps__n37;
wire sps__n38;
wire sps__n39;
wire sps__n40;
wire sps__n49;
wire sps__n52;
wire spc__n159;
wire sps__n54;
wire sps__n55;
wire sps__n57;
wire sps__n70;
wire sps__n71;
wire sps__n76;
wire sps__n77;
wire sps__n78;
wire sps__n79;
wire sps__n88;
wire sps__n89;
wire sps__n90;
wire sps__n97;
wire sps__n108;
wire sps__n109;
wire sps__n110;
wire sps__n117;
wire sps__n118;
wire sps__n119;
wire spc__n126;
wire spc__n127;
wire spc__n132;


OAI21_X1 i_0_0_181 (.ZN (n_119), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_28));
OAI21_X1 i_0_0_180 (.ZN (n_118), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_27));
OAI21_X1 i_0_0_179 (.ZN (n_117), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_28));
OAI21_X1 i_0_0_178 (.ZN (n_116), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_27));
OAI21_X1 i_0_0_177 (.ZN (n_115), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_26));
OAI21_X1 i_0_0_176 (.ZN (n_114), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_25));
OAI21_X1 i_0_0_175 (.ZN (n_113), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_26));
OAI21_X1 i_0_0_174 (.ZN (n_112), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_25));
OAI21_X1 i_0_0_173 (.ZN (n_111), .A (n_0_0_0), .B1 (n_0_0_45), .B2 (n_0_0_19));
OAI21_X1 i_0_0_172 (.ZN (n_110), .A (n_0_0_0), .B1 (n_0_0_45), .B2 (n_0_0_18));
OAI21_X1 i_0_0_171 (.ZN (n_109), .A (n_0_0_0), .B1 (n_0_0_44), .B2 (n_0_0_19));
OAI21_X1 i_0_0_170 (.ZN (n_108), .A (n_0_0_0), .B1 (n_0_0_44), .B2 (n_0_0_18));
OAI21_X1 i_0_0_169 (.ZN (n_107), .A (n_0_0_0), .B1 (n_0_0_45), .B2 (n_0_0_14));
OAI21_X1 i_0_0_168 (.ZN (n_106), .A (n_0_0_0), .B1 (n_0_0_45), .B2 (n_0_0_13));
NAND2_X1 i_0_0_167 (.ZN (n_0_0_45), .A1 (n_0_0_23), .A2 (n_0_0_41));
OAI21_X1 i_0_0_166 (.ZN (n_105), .A (n_0_0_0), .B1 (n_0_0_44), .B2 (n_0_0_14));
OAI21_X1 i_0_0_165 (.ZN (n_104), .A (n_0_0_0), .B1 (n_0_0_44), .B2 (n_0_0_13));
NAND2_X1 i_0_0_164 (.ZN (n_0_0_44), .A1 (n_0_0_21), .A2 (n_0_0_41));
OAI21_X1 i_0_0_163 (.ZN (n_103), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_19));
OAI21_X1 i_0_0_162 (.ZN (n_102), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_18));
OAI21_X1 i_0_0_161 (.ZN (n_101), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_19));
OAI21_X1 i_0_0_160 (.ZN (n_100), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_18));
OAI21_X1 i_0_0_159 (.ZN (n_99), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_14));
OAI21_X1 i_0_0_158 (.ZN (n_98), .A (n_0_0_0), .B1 (n_0_0_43), .B2 (n_0_0_13));
NAND2_X1 i_0_0_157 (.ZN (n_0_0_43), .A1 (n_0_0_16), .A2 (n_0_0_41));
OAI21_X1 i_0_0_156 (.ZN (n_97), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_14));
OAI21_X1 i_0_0_155 (.ZN (n_96), .A (n_0_0_0), .B1 (n_0_0_42), .B2 (n_0_0_13));
NAND2_X1 i_0_0_154 (.ZN (n_0_0_42), .A1 (n_0_0_7), .A2 (n_0_0_41));
NOR2_X1 i_0_0_153 (.ZN (n_0_0_41), .A1 (n_0_0_35), .A2 (n_0_0_29));
OAI21_X1 i_0_0_152 (.ZN (n_95), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_28));
OAI21_X1 i_0_0_151 (.ZN (n_94), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_27));
OAI21_X1 i_0_0_150 (.ZN (n_93), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_28));
OAI21_X1 i_0_0_149 (.ZN (n_92), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_27));
OAI21_X1 i_0_0_148 (.ZN (n_91), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_26));
OAI21_X1 i_0_0_147 (.ZN (n_90), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_25));
OAI21_X1 i_0_0_146 (.ZN (n_89), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_26));
OAI21_X1 i_0_0_145 (.ZN (n_88), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_25));
OAI21_X1 i_0_0_144 (.ZN (n_87), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_28));
OAI21_X1 i_0_0_143 (.ZN (n_86), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_27));
OAI21_X1 i_0_0_142 (.ZN (n_85), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_28));
OAI21_X1 i_0_0_141 (.ZN (n_84), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_27));
OAI21_X1 i_0_0_140 (.ZN (n_83), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_26));
OAI21_X1 i_0_0_139 (.ZN (n_82), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_25));
OAI21_X1 i_0_0_138 (.ZN (n_81), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_26));
OAI21_X1 i_0_0_137 (.ZN (n_80), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_25));
OAI21_X1 i_0_0_136 (.ZN (n_79), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_19));
OAI21_X1 i_0_0_135 (.ZN (n_78), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_18));
OAI21_X1 i_0_0_134 (.ZN (n_77), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_19));
OAI21_X1 i_0_0_133 (.ZN (n_76), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_18));
OAI21_X1 i_0_0_132 (.ZN (n_75), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_14));
OAI21_X1 i_0_0_131 (.ZN (n_74), .A (n_0_0_0), .B1 (n_0_0_40), .B2 (n_0_0_13));
NAND2_X1 i_0_0_130 (.ZN (n_0_0_40), .A1 (n_0_0_23), .A2 (n_0_0_36));
OAI21_X1 i_0_0_129 (.ZN (n_73), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_14));
OAI21_X1 i_0_0_128 (.ZN (n_72), .A (n_0_0_0), .B1 (n_0_0_39), .B2 (n_0_0_13));
NAND2_X1 i_0_0_127 (.ZN (n_0_0_39), .A1 (n_0_0_21), .A2 (n_0_0_36));
OAI21_X1 i_0_0_126 (.ZN (n_71), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_19));
OAI21_X1 i_0_0_125 (.ZN (n_70), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_18));
OAI21_X1 i_0_0_124 (.ZN (n_69), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_19));
OAI21_X1 i_0_0_123 (.ZN (n_68), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_18));
OAI21_X1 i_0_0_122 (.ZN (n_67), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_14));
OAI21_X1 i_0_0_121 (.ZN (n_66), .A (n_0_0_0), .B1 (n_0_0_38), .B2 (n_0_0_13));
NAND2_X1 i_0_0_120 (.ZN (n_0_0_38), .A1 (n_0_0_16), .A2 (n_0_0_36));
OAI21_X1 i_0_0_119 (.ZN (n_65), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_14));
OAI21_X1 i_0_0_118 (.ZN (n_64), .A (n_0_0_0), .B1 (n_0_0_37), .B2 (n_0_0_13));
NAND2_X1 i_0_0_117 (.ZN (n_0_0_37), .A1 (n_0_0_7), .A2 (n_0_0_36));
NOR2_X1 i_0_0_116 (.ZN (n_0_0_36), .A1 (n_0_0_35), .A2 (load_address[5]));
INV_X1 i_0_0_115 (.ZN (n_0_0_35), .A (load_address[6]));
OAI21_X1 i_0_0_114 (.ZN (n_63), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_28));
OAI21_X1 i_0_0_113 (.ZN (n_62), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_27));
OAI21_X1 i_0_0_112 (.ZN (n_61), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_28));
OAI21_X1 i_0_0_111 (.ZN (n_60), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_27));
OAI21_X1 i_0_0_110 (.ZN (n_59), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_26));
OAI21_X1 i_0_0_109 (.ZN (n_58), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_25));
OAI21_X1 i_0_0_108 (.ZN (n_57), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_26));
OAI21_X1 i_0_0_107 (.ZN (n_56), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_25));
OAI21_X1 i_0_0_106 (.ZN (n_55), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_28));
OAI21_X1 i_0_0_105 (.ZN (n_54), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_27));
OAI21_X1 i_0_0_104 (.ZN (n_53), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_28));
OAI21_X1 i_0_0_103 (.ZN (n_52), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_27));
OAI21_X1 i_0_0_102 (.ZN (n_51), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_26));
OAI21_X1 i_0_0_101 (.ZN (n_50), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_25));
OAI21_X1 i_0_0_100 (.ZN (n_49), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_26));
OAI21_X1 i_0_0_99 (.ZN (n_48), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_25));
OAI21_X1 i_0_0_98 (.ZN (n_47), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_19));
OAI21_X1 i_0_0_97 (.ZN (n_46), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_18));
OAI21_X1 i_0_0_96 (.ZN (n_45), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_19));
OAI21_X1 i_0_0_95 (.ZN (n_44), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_18));
OAI21_X1 i_0_0_94 (.ZN (n_43), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_14));
OAI21_X1 i_0_0_93 (.ZN (n_42), .A (n_0_0_0), .B1 (n_0_0_34), .B2 (n_0_0_13));
NAND2_X1 i_0_0_92 (.ZN (n_0_0_34), .A1 (n_0_0_23), .A2 (n_0_0_30));
OAI21_X1 i_0_0_91 (.ZN (n_41), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_14));
OAI21_X1 i_0_0_90 (.ZN (n_40), .A (n_0_0_0), .B1 (n_0_0_33), .B2 (n_0_0_13));
NAND2_X1 i_0_0_89 (.ZN (n_0_0_33), .A1 (n_0_0_21), .A2 (n_0_0_30));
OAI21_X1 i_0_0_88 (.ZN (n_39), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_19));
OAI21_X1 i_0_0_87 (.ZN (n_38), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_18));
OAI21_X1 i_0_0_86 (.ZN (n_37), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_19));
OAI21_X1 i_0_0_85 (.ZN (n_36), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_18));
OAI21_X1 i_0_0_84 (.ZN (n_35), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_14));
OAI21_X1 i_0_0_83 (.ZN (n_34), .A (n_0_0_0), .B1 (n_0_0_32), .B2 (n_0_0_13));
NAND2_X1 i_0_0_82 (.ZN (n_0_0_32), .A1 (n_0_0_16), .A2 (n_0_0_30));
OAI21_X1 i_0_0_81 (.ZN (n_33), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_14));
OAI21_X1 i_0_0_80 (.ZN (n_32), .A (n_0_0_0), .B1 (n_0_0_31), .B2 (n_0_0_13));
NAND2_X1 i_0_0_79 (.ZN (n_0_0_31), .A1 (n_0_0_7), .A2 (n_0_0_30));
NOR2_X1 i_0_0_78 (.ZN (n_0_0_30), .A1 (n_0_0_29), .A2 (load_address[6]));
INV_X1 i_0_0_77 (.ZN (n_0_0_29), .A (load_address[5]));
OAI21_X1 i_0_0_76 (.ZN (n_31), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_28));
OAI21_X1 i_0_0_75 (.ZN (n_30), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_27));
OAI21_X1 i_0_0_74 (.ZN (n_29), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_28));
OAI21_X1 i_0_0_73 (.ZN (n_28), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_27));
OAI21_X1 i_0_0_72 (.ZN (n_27), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_26));
OAI21_X1 i_0_0_71 (.ZN (n_26), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_25));
OAI21_X1 i_0_0_70 (.ZN (n_25), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_26));
OAI21_X1 i_0_0_69 (.ZN (n_24), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_25));
OAI21_X1 i_0_0_68 (.ZN (n_23), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_28));
OAI21_X1 i_0_0_67 (.ZN (n_22), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_27));
OAI21_X1 i_0_0_66 (.ZN (n_21), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_28));
NAND3_X1 i_0_0_65 (.ZN (n_0_0_28), .A1 (load_address[4]), .A2 (load_address[2]), .A3 (load_address[0]));
OAI21_X1 i_0_0_64 (.ZN (n_20), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_27));
NAND3_X1 i_0_0_63 (.ZN (n_0_0_27), .A1 (n_0_0_12), .A2 (load_address[4]), .A3 (load_address[2]));
OAI21_X1 i_0_0_62 (.ZN (n_19), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_26));
OAI21_X1 i_0_0_61 (.ZN (n_18), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_25));
OAI21_X1 i_0_0_60 (.ZN (n_17), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_26));
NAND3_X1 i_0_0_59 (.ZN (n_0_0_26), .A1 (n_0_0_11), .A2 (load_address[4]), .A3 (load_address[0]));
OAI21_X1 i_0_0_58 (.ZN (n_16), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_25));
NAND3_X1 i_0_0_57 (.ZN (n_0_0_25), .A1 (n_0_0_12), .A2 (n_0_0_11), .A3 (load_address[4]));
OAI21_X1 i_0_0_56 (.ZN (n_15), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_19));
OAI21_X1 i_0_0_55 (.ZN (n_14), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_18));
OAI21_X1 i_0_0_54 (.ZN (n_13), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_19));
OAI21_X1 i_0_0_53 (.ZN (n_12), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_18));
OAI21_X1 i_0_0_52 (.ZN (n_11), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_14));
OAI21_X1 i_0_0_51 (.ZN (n_10), .A (n_0_0_0), .B1 (n_0_0_24), .B2 (n_0_0_13));
NAND2_X1 i_0_0_50 (.ZN (n_0_0_24), .A1 (n_0_0_23), .A2 (n_0_0_8));
NOR2_X1 i_0_0_49 (.ZN (n_0_0_23), .A1 (n_0_0_15), .A2 (n_0_0_20));
OAI21_X1 i_0_0_48 (.ZN (n_9), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_14));
OAI21_X1 i_0_0_47 (.ZN (n_8), .A (n_0_0_0), .B1 (n_0_0_22), .B2 (n_0_0_13));
NAND2_X1 i_0_0_46 (.ZN (n_0_0_22), .A1 (n_0_0_21), .A2 (n_0_0_8));
NOR2_X1 i_0_0_45 (.ZN (n_0_0_21), .A1 (n_0_0_6), .A2 (n_0_0_20));
INV_X1 i_0_0_44 (.ZN (n_0_0_20), .A (load_address[3]));
OAI21_X1 i_0_0_43 (.ZN (n_7), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_19));
OAI21_X1 i_0_0_42 (.ZN (n_6), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_18));
OAI21_X1 i_0_0_41 (.ZN (n_5), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_19));
NAND3_X1 i_0_0_40 (.ZN (n_0_0_19), .A1 (n_0_0_10), .A2 (load_address[2]), .A3 (load_address[0]));
OAI21_X1 i_0_0_39 (.ZN (n_4), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_18));
NAND3_X1 i_0_0_38 (.ZN (n_0_0_18), .A1 (n_0_0_10), .A2 (n_0_0_12), .A3 (load_address[2]));
OAI21_X1 i_0_0_37 (.ZN (n_3), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_14));
OAI21_X1 i_0_0_36 (.ZN (n_2), .A (n_0_0_0), .B1 (n_0_0_17), .B2 (n_0_0_13));
NAND2_X1 i_0_0_35 (.ZN (n_0_0_17), .A1 (n_0_0_16), .A2 (n_0_0_8));
NOR2_X1 i_0_0_34 (.ZN (n_0_0_16), .A1 (n_0_0_15), .A2 (load_address[3]));
NAND2_X1 i_0_0_33 (.ZN (n_0_0_15), .A1 (n_0_0_4), .A2 (load_address[1]));
OAI21_X1 i_0_0_32 (.ZN (n_1), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_14));
NAND3_X1 i_0_0_31 (.ZN (n_0_0_14), .A1 (n_0_0_10), .A2 (n_0_0_11), .A3 (load_address[0]));
OAI21_X1 i_0_0_30 (.ZN (n_0), .A (n_0_0_0), .B1 (n_0_0_9), .B2 (n_0_0_13));
NAND3_X1 i_0_0_29 (.ZN (n_0_0_13), .A1 (n_0_0_10), .A2 (n_0_0_11), .A3 (n_0_0_12));
INV_X1 i_0_0_28 (.ZN (n_0_0_12), .A (load_address[0]));
INV_X1 i_0_0_27 (.ZN (n_0_0_11), .A (load_address[2]));
INV_X1 i_0_0_26 (.ZN (n_0_0_10), .A (load_address[4]));
NAND2_X1 i_0_0_25 (.ZN (n_0_0_9), .A1 (n_0_0_7), .A2 (n_0_0_8));
NOR2_X1 i_0_0_24 (.ZN (n_0_0_8), .A1 (load_address[6]), .A2 (load_address[5]));
NOR2_X1 i_0_0_23 (.ZN (n_0_0_7), .A1 (n_0_0_6), .A2 (load_address[3]));
NAND2_X1 i_0_0_22 (.ZN (n_0_0_6), .A1 (n_0_0_4), .A2 (n_0_0_5));
INV_X1 i_0_0_21 (.ZN (n_0_0_5), .A (load_address[1]));
AND4_X1 i_0_0_20 (.ZN (n_0_0_4), .A1 (n_0_0_1), .A2 (n_0_0_2), .A3 (n_0_0_3), .A4 (load_en));
INV_X1 i_0_0_19 (.ZN (n_0_0_3), .A (load_address[15]));
NOR4_X1 i_0_0_18 (.ZN (n_0_0_2), .A1 (load_address[10]), .A2 (load_address[9]), .A3 (load_address[8]), .A4 (load_address[7]));
NOR4_X1 i_0_0_17 (.ZN (n_0_0_1), .A1 (load_address[14]), .A2 (load_address[13]), .A3 (load_address[12]), .A4 (load_address[11]));
AND2_X1 i_0_0_16 (.ZN (\values[15] ), .A1 (n_0_0_0), .A2 (load_value[15]));
AND2_X1 i_0_0_15 (.ZN (\values[14] ), .A1 (n_0_0_0), .A2 (load_value[14]));
AND2_X1 i_0_0_14 (.ZN (\values[13] ), .A1 (n_0_0_0), .A2 (load_value[13]));
AND2_X1 i_0_0_13 (.ZN (\values[12] ), .A1 (n_0_0_0), .A2 (load_value[12]));
AND2_X1 i_0_0_12 (.ZN (\values[11] ), .A1 (n_0_0_0), .A2 (load_value[11]));
AND2_X1 i_0_0_11 (.ZN (\values[10] ), .A1 (n_0_0_0), .A2 (load_value[10]));
AND2_X1 i_0_0_10 (.ZN (\values[9] ), .A1 (n_0_0_0), .A2 (load_value[9]));
AND2_X1 i_0_0_9 (.ZN (\values[8] ), .A1 (n_0_0_0), .A2 (load_value[8]));
AND2_X4 i_0_0_8 (.ZN (\values[7] ), .A1 (n_0_0_0), .A2 (load_value[7]));
AND2_X1 i_0_0_7 (.ZN (\values[6] ), .A1 (n_0_0_0), .A2 (load_value[6]));
AND2_X4 i_0_0_6 (.ZN (\values[5] ), .A1 (n_0_0_0), .A2 (load_value[5]));
AND2_X1 i_0_0_5 (.ZN (\values[4] ), .A1 (n_0_0_0), .A2 (load_value[4]));
AND2_X1 i_0_0_4 (.ZN (\values[3] ), .A1 (n_0_0_0), .A2 (load_value[3]));
AND2_X4 i_0_0_3 (.ZN (\values[2] ), .A1 (n_0_0_0), .A2 (load_value[2]));
AND2_X1 i_0_0_2 (.ZN (\values[1] ), .A1 (n_0_0_0), .A2 (load_value[1]));
AND2_X1 i_0_0_1 (.ZN (\values[0] ), .A1 (n_0_0_0), .A2 (load_value[0]));
INV_X8 i_0_0_0 (.ZN (n_0_0_0), .A (reset));
DFF_X1 \values_reg[0][0]  (.Q (\values[0] [0] ), .CK (n_122_25), .D (sps__n5));
DFF_X1 \values_reg[0][1]  (.Q (\values[0] [1] ), .CK (n_122_25), .D (sps__n71));
DFF_X1 \values_reg[0][2]  (.Q (\values[0] [2] ), .CK (n_122_25), .D (spc__n159));
DFF_X1 \values_reg[0][3]  (.Q (\values[0] [3] ), .CK (n_122_25), .D (sps__n77));
DFF_X1 \values_reg[0][4]  (.Q (\values[0] [4] ), .CK (n_122_25), .D (sps__n90));
DFF_X1 \values_reg[0][5]  (.Q (\values[0] [5] ), .CK (n_122_25), .D (spc__n132));
DFF_X1 \values_reg[0][6]  (.Q (\values[0] [6] ), .CK (n_122_25), .D (sps__n117));
DFF_X1 \values_reg[0][7]  (.Q (\values[0] [7] ), .CK (n_122_25), .D (spc__n127));
DFF_X1 \values_reg[0][8]  (.Q (\values[0] [8] ), .CK (n_122_25), .D (sps__n97));
DFF_X1 \values_reg[0][9]  (.Q (\values[0] [9] ), .CK (n_122_25), .D (sps__n108));
DFF_X1 \values_reg[0][10]  (.Q (\values[0] [10] ), .CK (n_122_25), .D (sps__n1));
DFF_X1 \values_reg[0][11]  (.Q (\values[0] [11] ), .CK (n_122_25), .D (sps__n10));
DFF_X1 \values_reg[0][12]  (.Q (\values[0] [12] ), .CK (n_122_25), .D (sps__n57));
DFF_X1 \values_reg[0][13]  (.Q (\values[0] [13] ), .CK (n_122_25), .D (sps__n39));
DFF_X1 \values_reg[0][14]  (.Q (\values[0] [14] ), .CK (n_122_25), .D (sps__n27));
DFF_X1 \values_reg[0][15]  (.Q (\values[0] [15] ), .CK (n_122_25), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[0]_reg  (.GCK (n_122_25), .CK (clk), .E (n_0), .SE (1'b0 ));
DFF_X1 \values_reg[1][0]  (.Q (\values[1] [0] ), .CK (n_122_24), .D (sps__n5));
DFF_X1 \values_reg[1][1]  (.Q (\values[1] [1] ), .CK (n_122_24), .D (sps__n71));
DFF_X1 \values_reg[1][2]  (.Q (\values[1] [2] ), .CK (n_122_24), .D (spc__n159));
DFF_X1 \values_reg[1][3]  (.Q (\values[1] [3] ), .CK (n_122_24), .D (sps__n77));
DFF_X1 \values_reg[1][4]  (.Q (\values[1] [4] ), .CK (n_122_24), .D (sps__n89));
DFF_X1 \values_reg[1][5]  (.Q (\values[1] [5] ), .CK (n_122_24), .D (spc__n132));
DFF_X1 \values_reg[1][6]  (.Q (\values[1] [6] ), .CK (n_122_24), .D (sps__n117));
DFF_X1 \values_reg[1][7]  (.Q (\values[1] [7] ), .CK (n_122_24), .D (spc__n127));
DFF_X1 \values_reg[1][8]  (.Q (\values[1] [8] ), .CK (n_122_24), .D (sps__n97));
DFF_X1 \values_reg[1][9]  (.Q (\values[1] [9] ), .CK (n_122_24), .D (sps__n108));
DFF_X1 \values_reg[1][10]  (.Q (\values[1] [10] ), .CK (n_122_24), .D (sps__n1));
DFF_X1 \values_reg[1][11]  (.Q (\values[1] [11] ), .CK (n_122_24), .D (sps__n12));
DFF_X1 \values_reg[1][12]  (.Q (\values[1] [12] ), .CK (n_122_24), .D (sps__n54));
DFF_X1 \values_reg[1][13]  (.Q (\values[1] [13] ), .CK (n_122_24), .D (sps__n39));
DFF_X1 \values_reg[1][14]  (.Q (\values[1] [14] ), .CK (n_122_24), .D (sps__n27));
DFF_X1 \values_reg[1][15]  (.Q (\values[1] [15] ), .CK (n_122_24), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[1]_reg  (.GCK (n_122_24), .CK (clk), .E (n_1), .SE (1'b0 ));
DFF_X1 \values_reg[2][0]  (.Q (\values[2] [0] ), .CK (n_122_23), .D (sps__n5));
DFF_X1 \values_reg[2][1]  (.Q (\values[2] [1] ), .CK (n_122_23), .D (sps__n71));
DFF_X1 \values_reg[2][2]  (.Q (\values[2] [2] ), .CK (n_122_23), .D (spc__n159));
DFF_X1 \values_reg[2][3]  (.Q (\values[2] [3] ), .CK (n_122_23), .D (sps__n77));
DFF_X1 \values_reg[2][4]  (.Q (\values[2] [4] ), .CK (n_122_23), .D (sps__n89));
DFF_X1 \values_reg[2][5]  (.Q (\values[2] [5] ), .CK (n_122_23), .D (spc__n132));
DFF_X1 \values_reg[2][6]  (.Q (\values[2] [6] ), .CK (n_122_23), .D (sps__n118));
DFF_X1 \values_reg[2][7]  (.Q (\values[2] [7] ), .CK (n_122_23), .D (spc__n127));
DFF_X1 \values_reg[2][8]  (.Q (\values[2] [8] ), .CK (n_122_23), .D (sps__n97));
DFF_X1 \values_reg[2][9]  (.Q (\values[2] [9] ), .CK (n_122_23), .D (sps__n109));
DFF_X1 \values_reg[2][10]  (.Q (\values[2] [10] ), .CK (n_122_23), .D (sps__n1));
DFF_X1 \values_reg[2][11]  (.Q (\values[2] [11] ), .CK (n_122_23), .D (sps__n12));
DFF_X1 \values_reg[2][12]  (.Q (\values[2] [12] ), .CK (n_122_23), .D (sps__n54));
DFF_X1 \values_reg[2][13]  (.Q (\values[2] [13] ), .CK (n_122_23), .D (sps__n40));
DFF_X1 \values_reg[2][14]  (.Q (\values[2] [14] ), .CK (n_122_23), .D (sps__n28));
DFF_X1 \values_reg[2][15]  (.Q (\values[2] [15] ), .CK (n_122_23), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[2]_reg  (.GCK (n_122_23), .CK (clk), .E (n_2), .SE (1'b0 ));
DFF_X1 \values_reg[119][0]  (.Q (\values[119] [0] ), .CK (n_122_22), .D (sps__n5));
DFF_X1 \values_reg[119][1]  (.Q (\values[119] [1] ), .CK (n_122_22), .D (sps__n71));
DFF_X1 \values_reg[119][2]  (.Q (\values[119] [2] ), .CK (n_122_22), .D (spc__n157));
DFF_X1 \values_reg[119][3]  (.Q (\values[119] [3] ), .CK (n_122_22), .D (sps__n78));
DFF_X1 \values_reg[119][4]  (.Q (\values[119] [4] ), .CK (n_122_22), .D (sps__n89));
DFF_X1 \values_reg[119][5]  (.Q (\values[119] [5] ), .CK (n_122_22), .D (spc__n132));
DFF_X1 \values_reg[119][6]  (.Q (\values[119] [6] ), .CK (n_122_22), .D (sps__n118));
DFF_X1 \values_reg[119][7]  (.Q (\values[119] [7] ), .CK (n_122_22), .D (spc__n127));
DFF_X1 \values_reg[119][8]  (.Q (\values[119] [8] ), .CK (n_122_22), .D (sps__n97));
DFF_X1 \values_reg[119][9]  (.Q (\values[119] [9] ), .CK (n_122_22), .D (sps__n109));
DFF_X1 \values_reg[119][10]  (.Q (\values[119] [10] ), .CK (n_122_22), .D (sps__n1));
DFF_X1 \values_reg[119][11]  (.Q (\values[119] [11] ), .CK (n_122_22), .D (sps__n12));
DFF_X1 \values_reg[119][12]  (.Q (\values[119] [12] ), .CK (n_122_22), .D (sps__n52));
DFF_X1 \values_reg[119][13]  (.Q (\values[119] [13] ), .CK (n_122_22), .D (sps__n40));
DFF_X1 \values_reg[119][14]  (.Q (\values[119] [14] ), .CK (n_122_22), .D (sps__n28));
DFF_X1 \values_reg[119][15]  (.Q (\values[119] [15] ), .CK (n_122_22), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[119]_reg  (.GCK (n_122_22), .CK (clk), .E (n_119), .SE (1'b0 ));
DFF_X1 \values_reg[118][0]  (.Q (\values[118] [0] ), .CK (n_122_21), .D (sps__n5));
DFF_X1 \values_reg[118][1]  (.Q (\values[118] [1] ), .CK (n_122_21), .D (sps__n71));
DFF_X1 \values_reg[118][2]  (.Q (\values[118] [2] ), .CK (n_122_21), .D (spc__n159));
DFF_X1 \values_reg[118][3]  (.Q (\values[118] [3] ), .CK (n_122_21), .D (sps__n77));
DFF_X1 \values_reg[118][4]  (.Q (\values[118] [4] ), .CK (n_122_21), .D (sps__n90));
DFF_X1 \values_reg[118][5]  (.Q (\values[118] [5] ), .CK (n_122_21), .D (spc__n132));
DFF_X1 \values_reg[118][6]  (.Q (\values[118] [6] ), .CK (n_122_21), .D (sps__n118));
DFF_X1 \values_reg[118][7]  (.Q (\values[118] [7] ), .CK (n_122_21), .D (spc__n127));
DFF_X1 \values_reg[118][8]  (.Q (\values[118] [8] ), .CK (n_122_21), .D (sps__n97));
DFF_X1 \values_reg[118][9]  (.Q (\values[118] [9] ), .CK (n_122_21), .D (sps__n109));
DFF_X1 \values_reg[118][10]  (.Q (\values[118] [10] ), .CK (n_122_21), .D (sps__n1));
DFF_X1 \values_reg[118][11]  (.Q (\values[118] [11] ), .CK (n_122_21), .D (sps__n12));
DFF_X1 \values_reg[118][12]  (.Q (\values[118] [12] ), .CK (n_122_21), .D (sps__n54));
DFF_X1 \values_reg[118][13]  (.Q (\values[118] [13] ), .CK (n_122_21), .D (sps__n39));
DFF_X1 \values_reg[118][14]  (.Q (\values[118] [14] ), .CK (n_122_21), .D (sps__n27));
DFF_X1 \values_reg[118][15]  (.Q (\values[118] [15] ), .CK (n_122_21), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[118]_reg  (.GCK (n_122_21), .CK (clk), .E (n_118), .SE (1'b0 ));
DFF_X1 \values_reg[117][0]  (.Q (\values[117] [0] ), .CK (n_122_20), .D (sps__n5));
DFF_X1 \values_reg[117][1]  (.Q (\values[117] [1] ), .CK (n_122_20), .D (sps__n71));
DFF_X1 \values_reg[117][2]  (.Q (\values[117] [2] ), .CK (n_122_20), .D (spc__n157));
DFF_X1 \values_reg[117][3]  (.Q (\values[117] [3] ), .CK (n_122_20), .D (sps__n78));
DFF_X1 \values_reg[117][4]  (.Q (\values[117] [4] ), .CK (n_122_20), .D (sps__n89));
DFF_X1 \values_reg[117][5]  (.Q (\values[117] [5] ), .CK (n_122_20), .D (spc__n132));
DFF_X1 \values_reg[117][6]  (.Q (\values[117] [6] ), .CK (n_122_20), .D (sps__n118));
DFF_X1 \values_reg[117][7]  (.Q (\values[117] [7] ), .CK (n_122_20), .D (spc__n126));
DFF_X1 \values_reg[117][8]  (.Q (\values[117] [8] ), .CK (n_122_20), .D (sps__n97));
DFF_X1 \values_reg[117][9]  (.Q (\values[117] [9] ), .CK (n_122_20), .D (sps__n109));
DFF_X1 \values_reg[117][10]  (.Q (\values[117] [10] ), .CK (n_122_20), .D (sps__n1));
DFF_X1 \values_reg[117][11]  (.Q (\values[117] [11] ), .CK (n_122_20), .D (sps__n12));
DFF_X1 \values_reg[117][12]  (.Q (\values[117] [12] ), .CK (n_122_20), .D (sps__n55));
DFF_X1 \values_reg[117][13]  (.Q (\values[117] [13] ), .CK (n_122_20), .D (sps__n40));
DFF_X1 \values_reg[117][14]  (.Q (\values[117] [14] ), .CK (n_122_20), .D (sps__n28));
DFF_X1 \values_reg[117][15]  (.Q (\values[117] [15] ), .CK (n_122_20), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[117]_reg  (.GCK (n_122_20), .CK (clk), .E (n_117), .SE (1'b0 ));
DFF_X1 \values_reg[116][0]  (.Q (\values[116] [0] ), .CK (n_122_19), .D (sps__n5));
DFF_X1 \values_reg[116][1]  (.Q (\values[116] [1] ), .CK (n_122_19), .D (sps__n71));
DFF_X1 \values_reg[116][2]  (.Q (\values[116] [2] ), .CK (n_122_19), .D (spc__n157));
DFF_X1 \values_reg[116][3]  (.Q (\values[116] [3] ), .CK (n_122_19), .D (sps__n79));
DFF_X1 \values_reg[116][4]  (.Q (\values[116] [4] ), .CK (n_122_19), .D (sps__n89));
DFF_X1 \values_reg[116][5]  (.Q (\values[116] [5] ), .CK (n_122_19), .D (spc__n132));
DFF_X1 \values_reg[116][6]  (.Q (\values[116] [6] ), .CK (n_122_19), .D (sps__n118));
DFF_X1 \values_reg[116][7]  (.Q (\values[116] [7] ), .CK (n_122_19), .D (spc__n126));
DFF_X1 \values_reg[116][8]  (.Q (\values[116] [8] ), .CK (n_122_19), .D (sps__n97));
DFF_X1 \values_reg[116][9]  (.Q (\values[116] [9] ), .CK (n_122_19), .D (sps__n109));
DFF_X1 \values_reg[116][10]  (.Q (\values[116] [10] ), .CK (n_122_19), .D (sps__n1));
DFF_X1 \values_reg[116][11]  (.Q (\values[116] [11] ), .CK (n_122_19), .D (sps__n12));
DFF_X1 \values_reg[116][12]  (.Q (\values[116] [12] ), .CK (n_122_19), .D (sps__n55));
DFF_X1 \values_reg[116][13]  (.Q (\values[116] [13] ), .CK (n_122_19), .D (sps__n40));
DFF_X1 \values_reg[116][14]  (.Q (\values[116] [14] ), .CK (n_122_19), .D (sps__n28));
DFF_X1 \values_reg[116][15]  (.Q (\values[116] [15] ), .CK (n_122_19), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[116]_reg  (.GCK (n_122_19), .CK (clk), .E (n_116), .SE (1'b0 ));
DFF_X1 \values_reg[115][0]  (.Q (\values[115] [0] ), .CK (n_122_18), .D (sps__n5));
DFF_X1 \values_reg[115][1]  (.Q (\values[115] [1] ), .CK (n_122_18), .D (sps__n71));
DFF_X1 \values_reg[115][2]  (.Q (\values[115] [2] ), .CK (n_122_18), .D (spc__n159));
DFF_X1 \values_reg[115][3]  (.Q (\values[115] [3] ), .CK (n_122_18), .D (sps__n77));
DFF_X1 \values_reg[115][4]  (.Q (\values[115] [4] ), .CK (n_122_18), .D (sps__n90));
DFF_X1 \values_reg[115][5]  (.Q (\values[115] [5] ), .CK (n_122_18), .D (spc__n132));
DFF_X1 \values_reg[115][6]  (.Q (\values[115] [6] ), .CK (n_122_18), .D (sps__n117));
DFF_X1 \values_reg[115][7]  (.Q (\values[115] [7] ), .CK (n_122_18), .D (spc__n127));
DFF_X1 \values_reg[115][8]  (.Q (\values[115] [8] ), .CK (n_122_18), .D (sps__n97));
DFF_X1 \values_reg[115][9]  (.Q (\values[115] [9] ), .CK (n_122_18), .D (sps__n109));
DFF_X1 \values_reg[115][10]  (.Q (\values[115] [10] ), .CK (n_122_18), .D (sps__n1));
DFF_X1 \values_reg[115][11]  (.Q (\values[115] [11] ), .CK (n_122_18), .D (sps__n10));
DFF_X1 \values_reg[115][12]  (.Q (\values[115] [12] ), .CK (n_122_18), .D (sps__n54));
DFF_X1 \values_reg[115][13]  (.Q (\values[115] [13] ), .CK (n_122_18), .D (sps__n39));
DFF_X1 \values_reg[115][14]  (.Q (\values[115] [14] ), .CK (n_122_18), .D (sps__n27));
DFF_X1 \values_reg[115][15]  (.Q (\values[115] [15] ), .CK (n_122_18), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[115]_reg  (.GCK (n_122_18), .CK (clk), .E (n_115), .SE (1'b0 ));
DFF_X1 \values_reg[114][0]  (.Q (\values[114] [0] ), .CK (n_122_17), .D (sps__n5));
DFF_X1 \values_reg[114][1]  (.Q (\values[114] [1] ), .CK (n_122_17), .D (sps__n71));
DFF_X1 \values_reg[114][2]  (.Q (\values[114] [2] ), .CK (n_122_17), .D (spc__n159));
DFF_X1 \values_reg[114][3]  (.Q (\values[114] [3] ), .CK (n_122_17), .D (sps__n78));
DFF_X1 \values_reg[114][4]  (.Q (\values[114] [4] ), .CK (n_122_17), .D (sps__n90));
DFF_X1 \values_reg[114][5]  (.Q (\values[114] [5] ), .CK (n_122_17), .D (spc__n132));
DFF_X1 \values_reg[114][6]  (.Q (\values[114] [6] ), .CK (n_122_17), .D (sps__n117));
DFF_X1 \values_reg[114][7]  (.Q (\values[114] [7] ), .CK (n_122_17), .D (spc__n127));
DFF_X1 \values_reg[114][8]  (.Q (\values[114] [8] ), .CK (n_122_17), .D (sps__n97));
DFF_X1 \values_reg[114][9]  (.Q (\values[114] [9] ), .CK (n_122_17), .D (sps__n109));
DFF_X1 \values_reg[114][10]  (.Q (\values[114] [10] ), .CK (n_122_17), .D (sps__n1));
DFF_X1 \values_reg[114][11]  (.Q (\values[114] [11] ), .CK (n_122_17), .D (sps__n10));
DFF_X1 \values_reg[114][12]  (.Q (\values[114] [12] ), .CK (n_122_17), .D (sps__n52));
DFF_X1 \values_reg[114][13]  (.Q (\values[114] [13] ), .CK (n_122_17), .D (sps__n39));
DFF_X1 \values_reg[114][14]  (.Q (\values[114] [14] ), .CK (n_122_17), .D (sps__n27));
DFF_X1 \values_reg[114][15]  (.Q (\values[114] [15] ), .CK (n_122_17), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[114]_reg  (.GCK (n_122_17), .CK (clk), .E (n_114), .SE (1'b0 ));
DFF_X1 \values_reg[113][0]  (.Q (\values[113] [0] ), .CK (n_122_16), .D (sps__n5));
DFF_X1 \values_reg[113][1]  (.Q (\values[113] [1] ), .CK (n_122_16), .D (sps__n71));
DFF_X1 \values_reg[113][2]  (.Q (\values[113] [2] ), .CK (n_122_16), .D (spc__n157));
DFF_X1 \values_reg[113][3]  (.Q (\values[113] [3] ), .CK (n_122_16), .D (sps__n79));
DFF_X1 \values_reg[113][4]  (.Q (\values[113] [4] ), .CK (n_122_16), .D (sps__n89));
DFF_X1 \values_reg[113][5]  (.Q (\values[113] [5] ), .CK (n_122_16), .D (spc__n132));
DFF_X1 \values_reg[113][6]  (.Q (\values[113] [6] ), .CK (n_122_16), .D (sps__n118));
DFF_X1 \values_reg[113][7]  (.Q (\values[113] [7] ), .CK (n_122_16), .D (spc__n126));
DFF_X1 \values_reg[113][8]  (.Q (\values[113] [8] ), .CK (n_122_16), .D (sps__n97));
DFF_X1 \values_reg[113][9]  (.Q (\values[113] [9] ), .CK (n_122_16), .D (sps__n109));
DFF_X1 \values_reg[113][10]  (.Q (\values[113] [10] ), .CK (n_122_16), .D (sps__n1));
DFF_X1 \values_reg[113][11]  (.Q (\values[113] [11] ), .CK (n_122_16), .D (sps__n12));
DFF_X1 \values_reg[113][12]  (.Q (\values[113] [12] ), .CK (n_122_16), .D (sps__n55));
DFF_X1 \values_reg[113][13]  (.Q (\values[113] [13] ), .CK (n_122_16), .D (sps__n40));
DFF_X1 \values_reg[113][14]  (.Q (\values[113] [14] ), .CK (n_122_16), .D (sps__n28));
DFF_X1 \values_reg[113][15]  (.Q (\values[113] [15] ), .CK (n_122_16), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[113]_reg  (.GCK (n_122_16), .CK (clk), .E (n_113), .SE (1'b0 ));
DFF_X1 \values_reg[112][0]  (.Q (\values[112] [0] ), .CK (n_122_15), .D (sps__n5));
DFF_X1 \values_reg[112][1]  (.Q (\values[112] [1] ), .CK (n_122_15), .D (sps__n71));
DFF_X1 \values_reg[112][2]  (.Q (\values[112] [2] ), .CK (n_122_15), .D (spc__n157));
DFF_X1 \values_reg[112][3]  (.Q (\values[112] [3] ), .CK (n_122_15), .D (sps__n78));
DFF_X1 \values_reg[112][4]  (.Q (\values[112] [4] ), .CK (n_122_15), .D (sps__n89));
DFF_X1 \values_reg[112][5]  (.Q (\values[112] [5] ), .CK (n_122_15), .D (spc__n132));
DFF_X1 \values_reg[112][6]  (.Q (\values[112] [6] ), .CK (n_122_15), .D (sps__n118));
DFF_X1 \values_reg[112][7]  (.Q (\values[112] [7] ), .CK (n_122_15), .D (spc__n126));
DFF_X1 \values_reg[112][8]  (.Q (\values[112] [8] ), .CK (n_122_15), .D (sps__n97));
DFF_X1 \values_reg[112][9]  (.Q (\values[112] [9] ), .CK (n_122_15), .D (sps__n110));
DFF_X1 \values_reg[112][10]  (.Q (\values[112] [10] ), .CK (n_122_15), .D (sps__n1));
DFF_X1 \values_reg[112][11]  (.Q (\values[112] [11] ), .CK (n_122_15), .D (sps__n12));
DFF_X1 \values_reg[112][12]  (.Q (\values[112] [12] ), .CK (n_122_15), .D (sps__n55));
DFF_X1 \values_reg[112][13]  (.Q (\values[112] [13] ), .CK (n_122_15), .D (sps__n40));
DFF_X1 \values_reg[112][14]  (.Q (\values[112] [14] ), .CK (n_122_15), .D (sps__n28));
DFF_X1 \values_reg[112][15]  (.Q (\values[112] [15] ), .CK (n_122_15), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[112]_reg  (.GCK (n_122_15), .CK (clk), .E (n_112), .SE (1'b0 ));
DFF_X1 \values_reg[111][0]  (.Q (\values[111] [0] ), .CK (n_122_14), .D (sps__n5));
DFF_X1 \values_reg[111][1]  (.Q (\values[111] [1] ), .CK (n_122_14), .D (sps__n71));
DFF_X1 \values_reg[111][2]  (.Q (\values[111] [2] ), .CK (n_122_14), .D (spc__n159));
DFF_X1 \values_reg[111][3]  (.Q (\values[111] [3] ), .CK (n_122_14), .D (sps__n77));
DFF_X1 \values_reg[111][4]  (.Q (\values[111] [4] ), .CK (n_122_14), .D (sps__n90));
DFF_X1 \values_reg[111][5]  (.Q (\values[111] [5] ), .CK (n_122_14), .D (spc__n132));
DFF_X1 \values_reg[111][6]  (.Q (\values[111] [6] ), .CK (n_122_14), .D (sps__n117));
DFF_X1 \values_reg[111][7]  (.Q (\values[111] [7] ), .CK (n_122_14), .D (spc__n127));
DFF_X1 \values_reg[111][8]  (.Q (\values[111] [8] ), .CK (n_122_14), .D (sps__n97));
DFF_X1 \values_reg[111][9]  (.Q (\values[111] [9] ), .CK (n_122_14), .D (sps__n108));
DFF_X1 \values_reg[111][10]  (.Q (\values[111] [10] ), .CK (n_122_14), .D (sps__n1));
DFF_X1 \values_reg[111][11]  (.Q (\values[111] [11] ), .CK (n_122_14), .D (sps__n11));
DFF_X1 \values_reg[111][12]  (.Q (\values[111] [12] ), .CK (n_122_14), .D (sps__n57));
DFF_X1 \values_reg[111][13]  (.Q (\values[111] [13] ), .CK (n_122_14), .D (sps__n39));
DFF_X1 \values_reg[111][14]  (.Q (\values[111] [14] ), .CK (n_122_14), .D (sps__n25));
DFF_X1 \values_reg[111][15]  (.Q (\values[111] [15] ), .CK (n_122_14), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[111]_reg  (.GCK (n_122_14), .CK (clk), .E (n_111), .SE (1'b0 ));
DFF_X1 \values_reg[110][0]  (.Q (\values[110] [0] ), .CK (n_122_13), .D (sps__n5));
DFF_X1 \values_reg[110][1]  (.Q (\values[110] [1] ), .CK (n_122_13), .D (sps__n71));
DFF_X1 \values_reg[110][2]  (.Q (\values[110] [2] ), .CK (n_122_13), .D (spc__n159));
DFF_X1 \values_reg[110][3]  (.Q (\values[110] [3] ), .CK (n_122_13), .D (sps__n77));
DFF_X1 \values_reg[110][4]  (.Q (\values[110] [4] ), .CK (n_122_13), .D (sps__n90));
DFF_X1 \values_reg[110][5]  (.Q (\values[110] [5] ), .CK (n_122_13), .D (spc__n132));
DFF_X1 \values_reg[110][6]  (.Q (\values[110] [6] ), .CK (n_122_13), .D (sps__n117));
DFF_X1 \values_reg[110][7]  (.Q (\values[110] [7] ), .CK (n_122_13), .D (spc__n127));
DFF_X1 \values_reg[110][8]  (.Q (\values[110] [8] ), .CK (n_122_13), .D (sps__n97));
DFF_X1 \values_reg[110][9]  (.Q (\values[110] [9] ), .CK (n_122_13), .D (sps__n108));
DFF_X1 \values_reg[110][10]  (.Q (\values[110] [10] ), .CK (n_122_13), .D (sps__n1));
DFF_X1 \values_reg[110][11]  (.Q (\values[110] [11] ), .CK (n_122_13), .D (sps__n11));
DFF_X1 \values_reg[110][12]  (.Q (\values[110] [12] ), .CK (n_122_13), .D (sps__n57));
DFF_X1 \values_reg[110][13]  (.Q (\values[110] [13] ), .CK (n_122_13), .D (sps__n39));
DFF_X1 \values_reg[110][14]  (.Q (\values[110] [14] ), .CK (n_122_13), .D (sps__n25));
DFF_X1 \values_reg[110][15]  (.Q (\values[110] [15] ), .CK (n_122_13), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[110]_reg  (.GCK (n_122_13), .CK (clk), .E (n_110), .SE (1'b0 ));
DFF_X1 \values_reg[109][0]  (.Q (\values[109] [0] ), .CK (n_122_12), .D (sps__n5));
DFF_X1 \values_reg[109][1]  (.Q (\values[109] [1] ), .CK (n_122_12), .D (sps__n71));
DFF_X1 \values_reg[109][2]  (.Q (\values[109] [2] ), .CK (n_122_12), .D (spc__n158));
DFF_X1 \values_reg[109][3]  (.Q (\values[109] [3] ), .CK (n_122_12), .D (sps__n79));
DFF_X1 \values_reg[109][4]  (.Q (\values[109] [4] ), .CK (n_122_12), .D (sps__n89));
DFF_X1 \values_reg[109][5]  (.Q (\values[109] [5] ), .CK (n_122_12), .D (spc__n132));
DFF_X1 \values_reg[109][6]  (.Q (\values[109] [6] ), .CK (n_122_12), .D (sps__n119));
DFF_X1 \values_reg[109][7]  (.Q (\values[109] [7] ), .CK (n_122_12), .D (spc__n126));
DFF_X1 \values_reg[109][8]  (.Q (\values[109] [8] ), .CK (n_122_12), .D (sps__n97));
DFF_X1 \values_reg[109][9]  (.Q (\values[109] [9] ), .CK (n_122_12), .D (sps__n110));
DFF_X1 \values_reg[109][10]  (.Q (\values[109] [10] ), .CK (n_122_12), .D (sps__n1));
DFF_X1 \values_reg[109][11]  (.Q (\values[109] [11] ), .CK (n_122_12), .D (sps__n14));
DFF_X1 \values_reg[109][12]  (.Q (\values[109] [12] ), .CK (n_122_12), .D (sps__n52));
DFF_X1 \values_reg[109][13]  (.Q (\values[109] [13] ), .CK (n_122_12), .D (sps__n38));
DFF_X1 \values_reg[109][14]  (.Q (\values[109] [14] ), .CK (n_122_12), .D (sps__n28));
DFF_X1 \values_reg[109][15]  (.Q (\values[109] [15] ), .CK (n_122_12), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[109]_reg  (.GCK (n_122_12), .CK (clk), .E (n_109), .SE (1'b0 ));
DFF_X1 \values_reg[108][0]  (.Q (\values[108] [0] ), .CK (n_122_11), .D (sps__n5));
DFF_X1 \values_reg[108][1]  (.Q (\values[108] [1] ), .CK (n_122_11), .D (sps__n71));
DFF_X1 \values_reg[108][2]  (.Q (\values[108] [2] ), .CK (n_122_11), .D (spc__n157));
DFF_X1 \values_reg[108][3]  (.Q (\values[108] [3] ), .CK (n_122_11), .D (sps__n79));
DFF_X1 \values_reg[108][4]  (.Q (\values[108] [4] ), .CK (n_122_11), .D (sps__n89));
DFF_X1 \values_reg[108][5]  (.Q (\values[108] [5] ), .CK (n_122_11), .D (spc__n132));
DFF_X1 \values_reg[108][6]  (.Q (\values[108] [6] ), .CK (n_122_11), .D (sps__n119));
DFF_X1 \values_reg[108][7]  (.Q (\values[108] [7] ), .CK (n_122_11), .D (spc__n126));
DFF_X1 \values_reg[108][8]  (.Q (\values[108] [8] ), .CK (n_122_11), .D (sps__n97));
DFF_X1 \values_reg[108][9]  (.Q (\values[108] [9] ), .CK (n_122_11), .D (sps__n110));
DFF_X1 \values_reg[108][10]  (.Q (\values[108] [10] ), .CK (n_122_11), .D (sps__n1));
DFF_X1 \values_reg[108][11]  (.Q (\values[108] [11] ), .CK (n_122_11), .D (sps__n14));
DFF_X1 \values_reg[108][12]  (.Q (\values[108] [12] ), .CK (n_122_11), .D (sps__n52));
DFF_X1 \values_reg[108][13]  (.Q (\values[108] [13] ), .CK (n_122_11), .D (sps__n38));
DFF_X1 \values_reg[108][14]  (.Q (\values[108] [14] ), .CK (n_122_11), .D (sps__n28));
DFF_X1 \values_reg[108][15]  (.Q (\values[108] [15] ), .CK (n_122_11), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[108]_reg  (.GCK (n_122_11), .CK (clk), .E (n_108), .SE (1'b0 ));
DFF_X1 \values_reg[107][0]  (.Q (\values[107] [0] ), .CK (n_122_10), .D (sps__n5));
DFF_X1 \values_reg[107][1]  (.Q (\values[107] [1] ), .CK (n_122_10), .D (sps__n71));
DFF_X1 \values_reg[107][2]  (.Q (\values[107] [2] ), .CK (n_122_10), .D (spc__n159));
DFF_X1 \values_reg[107][3]  (.Q (\values[107] [3] ), .CK (n_122_10), .D (sps__n77));
DFF_X1 \values_reg[107][4]  (.Q (\values[107] [4] ), .CK (n_122_10), .D (sps__n90));
DFF_X1 \values_reg[107][5]  (.Q (\values[107] [5] ), .CK (n_122_10), .D (spc__n132));
DFF_X1 \values_reg[107][6]  (.Q (\values[107] [6] ), .CK (n_122_10), .D (sps__n117));
DFF_X1 \values_reg[107][7]  (.Q (\values[107] [7] ), .CK (n_122_10), .D (spc__n127));
DFF_X1 \values_reg[107][8]  (.Q (\values[107] [8] ), .CK (n_122_10), .D (sps__n97));
DFF_X1 \values_reg[107][9]  (.Q (\values[107] [9] ), .CK (n_122_10), .D (\values[9] ));
DFF_X1 \values_reg[107][10]  (.Q (\values[107] [10] ), .CK (n_122_10), .D (sps__n1));
DFF_X1 \values_reg[107][11]  (.Q (\values[107] [11] ), .CK (n_122_10), .D (sps__n11));
DFF_X1 \values_reg[107][12]  (.Q (\values[107] [12] ), .CK (n_122_10), .D (sps__n57));
DFF_X1 \values_reg[107][13]  (.Q (\values[107] [13] ), .CK (n_122_10), .D (sps__n39));
DFF_X1 \values_reg[107][14]  (.Q (\values[107] [14] ), .CK (n_122_10), .D (sps__n25));
DFF_X1 \values_reg[107][15]  (.Q (\values[107] [15] ), .CK (n_122_10), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[107]_reg  (.GCK (n_122_10), .CK (clk), .E (n_107), .SE (1'b0 ));
DFF_X1 \values_reg[106][0]  (.Q (\values[106] [0] ), .CK (n_122_9), .D (sps__n5));
DFF_X1 \values_reg[106][1]  (.Q (\values[106] [1] ), .CK (n_122_9), .D (sps__n71));
DFF_X1 \values_reg[106][2]  (.Q (\values[106] [2] ), .CK (n_122_9), .D (spc__n159));
DFF_X1 \values_reg[106][3]  (.Q (\values[106] [3] ), .CK (n_122_9), .D (sps__n76));
DFF_X1 \values_reg[106][4]  (.Q (\values[106] [4] ), .CK (n_122_9), .D (sps__n90));
DFF_X1 \values_reg[106][5]  (.Q (\values[106] [5] ), .CK (n_122_9), .D (spc__n132));
DFF_X1 \values_reg[106][6]  (.Q (\values[106] [6] ), .CK (n_122_9), .D (sps__n117));
DFF_X1 \values_reg[106][7]  (.Q (\values[106] [7] ), .CK (n_122_9), .D (spc__n127));
DFF_X1 \values_reg[106][8]  (.Q (\values[106] [8] ), .CK (n_122_9), .D (sps__n97));
DFF_X1 \values_reg[106][9]  (.Q (\values[106] [9] ), .CK (n_122_9), .D (sps__n108));
DFF_X1 \values_reg[106][10]  (.Q (\values[106] [10] ), .CK (n_122_9), .D (sps__n1));
DFF_X1 \values_reg[106][11]  (.Q (\values[106] [11] ), .CK (n_122_9), .D (sps__n10));
DFF_X1 \values_reg[106][12]  (.Q (\values[106] [12] ), .CK (n_122_9), .D (sps__n57));
DFF_X1 \values_reg[106][13]  (.Q (\values[106] [13] ), .CK (n_122_9), .D (sps__n37));
DFF_X1 \values_reg[106][14]  (.Q (\values[106] [14] ), .CK (n_122_9), .D (sps__n25));
DFF_X1 \values_reg[106][15]  (.Q (\values[106] [15] ), .CK (n_122_9), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[106]_reg  (.GCK (n_122_9), .CK (clk), .E (n_106), .SE (1'b0 ));
DFF_X1 \values_reg[105][0]  (.Q (\values[105] [0] ), .CK (n_122_8), .D (sps__n5));
DFF_X1 \values_reg[105][1]  (.Q (\values[105] [1] ), .CK (n_122_8), .D (sps__n71));
DFF_X1 \values_reg[105][2]  (.Q (\values[105] [2] ), .CK (n_122_8), .D (spc__n158));
DFF_X1 \values_reg[105][3]  (.Q (\values[105] [3] ), .CK (n_122_8), .D (sps__n77));
DFF_X1 \values_reg[105][4]  (.Q (\values[105] [4] ), .CK (n_122_8), .D (sps__n90));
DFF_X1 \values_reg[105][5]  (.Q (\values[105] [5] ), .CK (n_122_8), .D (spc__n132));
DFF_X1 \values_reg[105][6]  (.Q (\values[105] [6] ), .CK (n_122_8), .D (sps__n119));
DFF_X1 \values_reg[105][7]  (.Q (\values[105] [7] ), .CK (n_122_8), .D (spc__n126));
DFF_X1 \values_reg[105][8]  (.Q (\values[105] [8] ), .CK (n_122_8), .D (sps__n97));
DFF_X1 \values_reg[105][9]  (.Q (\values[105] [9] ), .CK (n_122_8), .D (sps__n110));
DFF_X1 \values_reg[105][10]  (.Q (\values[105] [10] ), .CK (n_122_8), .D (sps__n1));
DFF_X1 \values_reg[105][11]  (.Q (\values[105] [11] ), .CK (n_122_8), .D (sps__n14));
DFF_X1 \values_reg[105][12]  (.Q (\values[105] [12] ), .CK (n_122_8), .D (sps__n52));
DFF_X1 \values_reg[105][13]  (.Q (\values[105] [13] ), .CK (n_122_8), .D (sps__n38));
DFF_X1 \values_reg[105][14]  (.Q (\values[105] [14] ), .CK (n_122_8), .D (sps__n25));
DFF_X1 \values_reg[105][15]  (.Q (\values[105] [15] ), .CK (n_122_8), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[105]_reg  (.GCK (n_122_8), .CK (clk), .E (n_105), .SE (1'b0 ));
DFF_X1 \values_reg[104][0]  (.Q (\values[104] [0] ), .CK (n_122_7), .D (sps__n5));
DFF_X1 \values_reg[104][1]  (.Q (\values[104] [1] ), .CK (n_122_7), .D (sps__n71));
DFF_X1 \values_reg[104][2]  (.Q (\values[104] [2] ), .CK (n_122_7), .D (spc__n158));
DFF_X1 \values_reg[104][3]  (.Q (\values[104] [3] ), .CK (n_122_7), .D (sps__n77));
DFF_X1 \values_reg[104][4]  (.Q (\values[104] [4] ), .CK (n_122_7), .D (sps__n90));
DFF_X1 \values_reg[104][5]  (.Q (\values[104] [5] ), .CK (n_122_7), .D (spc__n132));
DFF_X1 \values_reg[104][6]  (.Q (\values[104] [6] ), .CK (n_122_7), .D (sps__n119));
DFF_X1 \values_reg[104][7]  (.Q (\values[104] [7] ), .CK (n_122_7), .D (spc__n126));
DFF_X1 \values_reg[104][8]  (.Q (\values[104] [8] ), .CK (n_122_7), .D (sps__n97));
DFF_X1 \values_reg[104][9]  (.Q (\values[104] [9] ), .CK (n_122_7), .D (\values[9] ));
DFF_X1 \values_reg[104][10]  (.Q (\values[104] [10] ), .CK (n_122_7), .D (sps__n1));
DFF_X1 \values_reg[104][11]  (.Q (\values[104] [11] ), .CK (n_122_7), .D (sps__n10));
DFF_X1 \values_reg[104][12]  (.Q (\values[104] [12] ), .CK (n_122_7), .D (sps__n52));
DFF_X1 \values_reg[104][13]  (.Q (\values[104] [13] ), .CK (n_122_7), .D (sps__n38));
DFF_X1 \values_reg[104][14]  (.Q (\values[104] [14] ), .CK (n_122_7), .D (sps__n28));
DFF_X1 \values_reg[104][15]  (.Q (\values[104] [15] ), .CK (n_122_7), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[104]_reg  (.GCK (n_122_7), .CK (clk), .E (n_104), .SE (1'b0 ));
DFF_X1 \values_reg[103][0]  (.Q (\values[103] [0] ), .CK (n_122_6), .D (sps__n5));
DFF_X1 \values_reg[103][1]  (.Q (\values[103] [1] ), .CK (n_122_6), .D (sps__n71));
DFF_X1 \values_reg[103][2]  (.Q (\values[103] [2] ), .CK (n_122_6), .D (spc__n159));
DFF_X1 \values_reg[103][3]  (.Q (\values[103] [3] ), .CK (n_122_6), .D (sps__n77));
DFF_X1 \values_reg[103][4]  (.Q (\values[103] [4] ), .CK (n_122_6), .D (sps__n90));
DFF_X1 \values_reg[103][5]  (.Q (\values[103] [5] ), .CK (n_122_6), .D (spc__n132));
DFF_X1 \values_reg[103][6]  (.Q (\values[103] [6] ), .CK (n_122_6), .D (sps__n117));
DFF_X1 \values_reg[103][7]  (.Q (\values[103] [7] ), .CK (n_122_6), .D (spc__n127));
DFF_X1 \values_reg[103][8]  (.Q (\values[103] [8] ), .CK (n_122_6), .D (sps__n97));
DFF_X1 \values_reg[103][9]  (.Q (\values[103] [9] ), .CK (n_122_6), .D (sps__n108));
DFF_X1 \values_reg[103][10]  (.Q (\values[103] [10] ), .CK (n_122_6), .D (sps__n1));
DFF_X1 \values_reg[103][11]  (.Q (\values[103] [11] ), .CK (n_122_6), .D (sps__n10));
DFF_X1 \values_reg[103][12]  (.Q (\values[103] [12] ), .CK (n_122_6), .D (sps__n52));
DFF_X1 \values_reg[103][13]  (.Q (\values[103] [13] ), .CK (n_122_6), .D (sps__n39));
DFF_X1 \values_reg[103][14]  (.Q (\values[103] [14] ), .CK (n_122_6), .D (sps__n27));
DFF_X1 \values_reg[103][15]  (.Q (\values[103] [15] ), .CK (n_122_6), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[103]_reg  (.GCK (n_122_6), .CK (clk), .E (n_103), .SE (1'b0 ));
DFF_X1 \values_reg[102][0]  (.Q (\values[102] [0] ), .CK (n_122_5), .D (sps__n5));
DFF_X1 \values_reg[102][1]  (.Q (\values[102] [1] ), .CK (n_122_5), .D (sps__n71));
DFF_X1 \values_reg[102][2]  (.Q (\values[102] [2] ), .CK (n_122_5), .D (\values[2] ));
DFF_X1 \values_reg[102][3]  (.Q (\values[102] [3] ), .CK (n_122_5), .D (sps__n77));
DFF_X1 \values_reg[102][4]  (.Q (\values[102] [4] ), .CK (n_122_5), .D (sps__n90));
DFF_X1 \values_reg[102][5]  (.Q (\values[102] [5] ), .CK (n_122_5), .D (spc__n132));
DFF_X1 \values_reg[102][6]  (.Q (\values[102] [6] ), .CK (n_122_5), .D (\values[6] ));
DFF_X1 \values_reg[102][7]  (.Q (\values[102] [7] ), .CK (n_122_5), .D (spc__n127));
DFF_X1 \values_reg[102][8]  (.Q (\values[102] [8] ), .CK (n_122_5), .D (sps__n97));
DFF_X1 \values_reg[102][9]  (.Q (\values[102] [9] ), .CK (n_122_5), .D (sps__n108));
DFF_X1 \values_reg[102][10]  (.Q (\values[102] [10] ), .CK (n_122_5), .D (sps__n1));
DFF_X1 \values_reg[102][11]  (.Q (\values[102] [11] ), .CK (n_122_5), .D (sps__n10));
DFF_X1 \values_reg[102][12]  (.Q (\values[102] [12] ), .CK (n_122_5), .D (sps__n52));
DFF_X1 \values_reg[102][13]  (.Q (\values[102] [13] ), .CK (n_122_5), .D (sps__n39));
DFF_X1 \values_reg[102][14]  (.Q (\values[102] [14] ), .CK (n_122_5), .D (sps__n28));
DFF_X1 \values_reg[102][15]  (.Q (\values[102] [15] ), .CK (n_122_5), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[102]_reg  (.GCK (n_122_5), .CK (clk), .E (n_102), .SE (1'b0 ));
DFF_X1 \values_reg[101][0]  (.Q (\values[101] [0] ), .CK (n_122_4), .D (sps__n5));
DFF_X1 \values_reg[101][1]  (.Q (\values[101] [1] ), .CK (n_122_4), .D (sps__n71));
DFF_X1 \values_reg[101][2]  (.Q (\values[101] [2] ), .CK (n_122_4), .D (spc__n157));
DFF_X1 \values_reg[101][3]  (.Q (\values[101] [3] ), .CK (n_122_4), .D (sps__n76));
DFF_X1 \values_reg[101][4]  (.Q (\values[101] [4] ), .CK (n_122_4), .D (sps__n88));
DFF_X1 \values_reg[101][5]  (.Q (\values[101] [5] ), .CK (n_122_4), .D (spc__n132));
DFF_X1 \values_reg[101][6]  (.Q (\values[101] [6] ), .CK (n_122_4), .D (\values[6] ));
DFF_X1 \values_reg[101][7]  (.Q (\values[101] [7] ), .CK (n_122_4), .D (\values[7] ));
DFF_X1 \values_reg[101][8]  (.Q (\values[101] [8] ), .CK (n_122_4), .D (sps__n97));
DFF_X1 \values_reg[101][9]  (.Q (\values[101] [9] ), .CK (n_122_4), .D (sps__n110));
DFF_X1 \values_reg[101][10]  (.Q (\values[101] [10] ), .CK (n_122_4), .D (sps__n1));
DFF_X1 \values_reg[101][11]  (.Q (\values[101] [11] ), .CK (n_122_4), .D (sps__n10));
DFF_X1 \values_reg[101][12]  (.Q (\values[101] [12] ), .CK (n_122_4), .D (sps__n52));
DFF_X1 \values_reg[101][13]  (.Q (\values[101] [13] ), .CK (n_122_4), .D (sps__n37));
DFF_X1 \values_reg[101][14]  (.Q (\values[101] [14] ), .CK (n_122_4), .D (sps__n28));
DFF_X1 \values_reg[101][15]  (.Q (\values[101] [15] ), .CK (n_122_4), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[101]_reg  (.GCK (n_122_4), .CK (clk), .E (n_101), .SE (1'b0 ));
DFF_X1 \values_reg[100][0]  (.Q (\values[100] [0] ), .CK (n_122_3), .D (sps__n5));
DFF_X1 \values_reg[100][1]  (.Q (\values[100] [1] ), .CK (n_122_3), .D (sps__n71));
DFF_X1 \values_reg[100][2]  (.Q (\values[100] [2] ), .CK (n_122_3), .D (spc__n157));
DFF_X1 \values_reg[100][3]  (.Q (\values[100] [3] ), .CK (n_122_3), .D (sps__n78));
DFF_X1 \values_reg[100][4]  (.Q (\values[100] [4] ), .CK (n_122_3), .D (sps__n89));
DFF_X1 \values_reg[100][5]  (.Q (\values[100] [5] ), .CK (n_122_3), .D (spc__n132));
DFF_X1 \values_reg[100][6]  (.Q (\values[100] [6] ), .CK (n_122_3), .D (sps__n118));
DFF_X1 \values_reg[100][7]  (.Q (\values[100] [7] ), .CK (n_122_3), .D (\values[7] ));
DFF_X1 \values_reg[100][8]  (.Q (\values[100] [8] ), .CK (n_122_3), .D (sps__n97));
DFF_X1 \values_reg[100][9]  (.Q (\values[100] [9] ), .CK (n_122_3), .D (sps__n110));
DFF_X1 \values_reg[100][10]  (.Q (\values[100] [10] ), .CK (n_122_3), .D (sps__n1));
DFF_X1 \values_reg[100][11]  (.Q (\values[100] [11] ), .CK (n_122_3), .D (sps__n12));
DFF_X1 \values_reg[100][12]  (.Q (\values[100] [12] ), .CK (n_122_3), .D (sps__n52));
DFF_X1 \values_reg[100][13]  (.Q (\values[100] [13] ), .CK (n_122_3), .D (sps__n37));
DFF_X1 \values_reg[100][14]  (.Q (\values[100] [14] ), .CK (n_122_3), .D (sps__n28));
DFF_X1 \values_reg[100][15]  (.Q (\values[100] [15] ), .CK (n_122_3), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[100]_reg  (.GCK (n_122_3), .CK (clk), .E (n_100), .SE (1'b0 ));
DFF_X1 \values_reg[99][0]  (.Q (\values[99] [0] ), .CK (n_122_2), .D (sps__n5));
DFF_X1 \values_reg[99][1]  (.Q (\values[99] [1] ), .CK (n_122_2), .D (sps__n71));
DFF_X1 \values_reg[99][2]  (.Q (\values[99] [2] ), .CK (n_122_2), .D (spc__n157));
DFF_X1 \values_reg[99][3]  (.Q (\values[99] [3] ), .CK (n_122_2), .D (sps__n78));
DFF_X1 \values_reg[99][4]  (.Q (\values[99] [4] ), .CK (n_122_2), .D (sps__n89));
DFF_X1 \values_reg[99][5]  (.Q (\values[99] [5] ), .CK (n_122_2), .D (spc__n132));
DFF_X1 \values_reg[99][6]  (.Q (\values[99] [6] ), .CK (n_122_2), .D (sps__n118));
DFF_X1 \values_reg[99][7]  (.Q (\values[99] [7] ), .CK (n_122_2), .D (spc__n126));
DFF_X1 \values_reg[99][8]  (.Q (\values[99] [8] ), .CK (n_122_2), .D (sps__n97));
DFF_X1 \values_reg[99][9]  (.Q (\values[99] [9] ), .CK (n_122_2), .D (sps__n109));
DFF_X1 \values_reg[99][10]  (.Q (\values[99] [10] ), .CK (n_122_2), .D (sps__n1));
DFF_X1 \values_reg[99][11]  (.Q (\values[99] [11] ), .CK (n_122_2), .D (sps__n12));
DFF_X1 \values_reg[99][12]  (.Q (\values[99] [12] ), .CK (n_122_2), .D (sps__n55));
DFF_X1 \values_reg[99][13]  (.Q (\values[99] [13] ), .CK (n_122_2), .D (sps__n40));
DFF_X1 \values_reg[99][14]  (.Q (\values[99] [14] ), .CK (n_122_2), .D (sps__n28));
DFF_X1 \values_reg[99][15]  (.Q (\values[99] [15] ), .CK (n_122_2), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[99]_reg  (.GCK (n_122_2), .CK (clk), .E (n_99), .SE (1'b0 ));
DFF_X1 \values_reg[98][0]  (.Q (\values[98] [0] ), .CK (n_122_1), .D (sps__n5));
DFF_X1 \values_reg[98][1]  (.Q (\values[98] [1] ), .CK (n_122_1), .D (sps__n71));
DFF_X1 \values_reg[98][2]  (.Q (\values[98] [2] ), .CK (n_122_1), .D (spc__n159));
DFF_X1 \values_reg[98][3]  (.Q (\values[98] [3] ), .CK (n_122_1), .D (sps__n78));
DFF_X1 \values_reg[98][4]  (.Q (\values[98] [4] ), .CK (n_122_1), .D (sps__n89));
DFF_X1 \values_reg[98][5]  (.Q (\values[98] [5] ), .CK (n_122_1), .D (spc__n132));
DFF_X1 \values_reg[98][6]  (.Q (\values[98] [6] ), .CK (n_122_1), .D (sps__n118));
DFF_X1 \values_reg[98][7]  (.Q (\values[98] [7] ), .CK (n_122_1), .D (spc__n126));
DFF_X1 \values_reg[98][8]  (.Q (\values[98] [8] ), .CK (n_122_1), .D (sps__n97));
DFF_X1 \values_reg[98][9]  (.Q (\values[98] [9] ), .CK (n_122_1), .D (sps__n109));
DFF_X1 \values_reg[98][10]  (.Q (\values[98] [10] ), .CK (n_122_1), .D (sps__n1));
DFF_X1 \values_reg[98][11]  (.Q (\values[98] [11] ), .CK (n_122_1), .D (sps__n12));
DFF_X1 \values_reg[98][12]  (.Q (\values[98] [12] ), .CK (n_122_1), .D (sps__n54));
DFF_X1 \values_reg[98][13]  (.Q (\values[98] [13] ), .CK (n_122_1), .D (sps__n40));
DFF_X1 \values_reg[98][14]  (.Q (\values[98] [14] ), .CK (n_122_1), .D (sps__n28));
DFF_X1 \values_reg[98][15]  (.Q (\values[98] [15] ), .CK (n_122_1), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[98]_reg  (.GCK (n_122_1), .CK (clk), .E (n_98), .SE (1'b0 ));
DFF_X1 \values_reg[97][0]  (.Q (\values[97] [0] ), .CK (n_122_0), .D (sps__n5));
DFF_X1 \values_reg[97][1]  (.Q (\values[97] [1] ), .CK (n_122_0), .D (sps__n71));
DFF_X1 \values_reg[97][2]  (.Q (\values[97] [2] ), .CK (n_122_0), .D (spc__n157));
DFF_X1 \values_reg[97][3]  (.Q (\values[97] [3] ), .CK (n_122_0), .D (sps__n79));
DFF_X1 \values_reg[97][4]  (.Q (\values[97] [4] ), .CK (n_122_0), .D (sps__n89));
DFF_X1 \values_reg[97][5]  (.Q (\values[97] [5] ), .CK (n_122_0), .D (spc__n132));
DFF_X1 \values_reg[97][6]  (.Q (\values[97] [6] ), .CK (n_122_0), .D (sps__n118));
DFF_X1 \values_reg[97][7]  (.Q (\values[97] [7] ), .CK (n_122_0), .D (spc__n126));
DFF_X1 \values_reg[97][8]  (.Q (\values[97] [8] ), .CK (n_122_0), .D (sps__n97));
DFF_X1 \values_reg[97][9]  (.Q (\values[97] [9] ), .CK (n_122_0), .D (sps__n109));
DFF_X1 \values_reg[97][10]  (.Q (\values[97] [10] ), .CK (n_122_0), .D (sps__n1));
DFF_X1 \values_reg[97][11]  (.Q (\values[97] [11] ), .CK (n_122_0), .D (sps__n12));
DFF_X1 \values_reg[97][12]  (.Q (\values[97] [12] ), .CK (n_122_0), .D (sps__n55));
DFF_X1 \values_reg[97][13]  (.Q (\values[97] [13] ), .CK (n_122_0), .D (sps__n40));
DFF_X1 \values_reg[97][14]  (.Q (\values[97] [14] ), .CK (n_122_0), .D (sps__n28));
DFF_X1 \values_reg[97][15]  (.Q (\values[97] [15] ), .CK (n_122_0), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[97]_reg  (.GCK (n_122_0), .CK (clk), .E (n_97), .SE (1'b0 ));
DFF_X1 \values_reg[26][0]  (.Q (\values[26] [0] ), .CK (n_121_93), .D (sps__n5));
DFF_X1 \values_reg[26][1]  (.Q (\values[26] [1] ), .CK (n_121_93), .D (sps__n71));
DFF_X1 \values_reg[26][2]  (.Q (\values[26] [2] ), .CK (n_121_93), .D (spc__n159));
DFF_X1 \values_reg[26][3]  (.Q (\values[26] [3] ), .CK (n_121_93), .D (sps__n77));
DFF_X1 \values_reg[26][4]  (.Q (\values[26] [4] ), .CK (n_121_93), .D (sps__n90));
DFF_X1 \values_reg[26][5]  (.Q (\values[26] [5] ), .CK (n_121_93), .D (spc__n132));
DFF_X1 \values_reg[26][6]  (.Q (\values[26] [6] ), .CK (n_121_93), .D (sps__n117));
DFF_X1 \values_reg[26][7]  (.Q (\values[26] [7] ), .CK (n_121_93), .D (spc__n127));
DFF_X1 \values_reg[26][8]  (.Q (\values[26] [8] ), .CK (n_121_93), .D (sps__n97));
DFF_X1 \values_reg[26][9]  (.Q (\values[26] [9] ), .CK (n_121_93), .D (sps__n108));
DFF_X1 \values_reg[26][10]  (.Q (\values[26] [10] ), .CK (n_121_93), .D (sps__n1));
DFF_X1 \values_reg[26][11]  (.Q (\values[26] [11] ), .CK (n_121_93), .D (sps__n11));
DFF_X1 \values_reg[26][12]  (.Q (\values[26] [12] ), .CK (n_121_93), .D (sps__n57));
DFF_X1 \values_reg[26][13]  (.Q (\values[26] [13] ), .CK (n_121_93), .D (sps__n39));
DFF_X1 \values_reg[26][14]  (.Q (\values[26] [14] ), .CK (n_121_93), .D (sps__n28));
DFF_X1 \values_reg[26][15]  (.Q (\values[26] [15] ), .CK (n_121_93), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[26]_reg  (.GCK (n_121_93), .CK (clk), .E (n_26), .SE (1'b0 ));
DFF_X1 \values_reg[27][0]  (.Q (\values[27] [0] ), .CK (n_121_92), .D (sps__n5));
DFF_X1 \values_reg[27][1]  (.Q (\values[27] [1] ), .CK (n_121_92), .D (sps__n71));
DFF_X1 \values_reg[27][2]  (.Q (\values[27] [2] ), .CK (n_121_92), .D (spc__n159));
DFF_X1 \values_reg[27][3]  (.Q (\values[27] [3] ), .CK (n_121_92), .D (sps__n77));
DFF_X1 \values_reg[27][4]  (.Q (\values[27] [4] ), .CK (n_121_92), .D (sps__n90));
DFF_X1 \values_reg[27][5]  (.Q (\values[27] [5] ), .CK (n_121_92), .D (spc__n132));
DFF_X1 \values_reg[27][6]  (.Q (\values[27] [6] ), .CK (n_121_92), .D (sps__n117));
DFF_X1 \values_reg[27][7]  (.Q (\values[27] [7] ), .CK (n_121_92), .D (spc__n127));
DFF_X1 \values_reg[27][8]  (.Q (\values[27] [8] ), .CK (n_121_92), .D (sps__n97));
DFF_X1 \values_reg[27][9]  (.Q (\values[27] [9] ), .CK (n_121_92), .D (sps__n108));
DFF_X1 \values_reg[27][10]  (.Q (\values[27] [10] ), .CK (n_121_92), .D (sps__n1));
DFF_X1 \values_reg[27][11]  (.Q (\values[27] [11] ), .CK (n_121_92), .D (sps__n11));
DFF_X1 \values_reg[27][12]  (.Q (\values[27] [12] ), .CK (n_121_92), .D (sps__n57));
DFF_X1 \values_reg[27][13]  (.Q (\values[27] [13] ), .CK (n_121_92), .D (sps__n39));
DFF_X1 \values_reg[27][14]  (.Q (\values[27] [14] ), .CK (n_121_92), .D (sps__n28));
DFF_X1 \values_reg[27][15]  (.Q (\values[27] [15] ), .CK (n_121_92), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[27]_reg  (.GCK (n_121_92), .CK (clk), .E (n_27), .SE (1'b0 ));
DFF_X1 \values_reg[28][0]  (.Q (\values[28] [0] ), .CK (n_121_91), .D (sps__n5));
DFF_X1 \values_reg[28][1]  (.Q (\values[28] [1] ), .CK (n_121_91), .D (sps__n71));
DFF_X1 \values_reg[28][2]  (.Q (\values[28] [2] ), .CK (n_121_91), .D (spc__n159));
DFF_X1 \values_reg[28][3]  (.Q (\values[28] [3] ), .CK (n_121_91), .D (sps__n77));
DFF_X1 \values_reg[28][4]  (.Q (\values[28] [4] ), .CK (n_121_91), .D (sps__n89));
DFF_X1 \values_reg[28][5]  (.Q (\values[28] [5] ), .CK (n_121_91), .D (spc__n132));
DFF_X1 \values_reg[28][6]  (.Q (\values[28] [6] ), .CK (n_121_91), .D (sps__n117));
DFF_X1 \values_reg[28][7]  (.Q (\values[28] [7] ), .CK (n_121_91), .D (spc__n127));
DFF_X1 \values_reg[28][8]  (.Q (\values[28] [8] ), .CK (n_121_91), .D (sps__n97));
DFF_X1 \values_reg[28][9]  (.Q (\values[28] [9] ), .CK (n_121_91), .D (sps__n109));
DFF_X1 \values_reg[28][10]  (.Q (\values[28] [10] ), .CK (n_121_91), .D (sps__n1));
DFF_X1 \values_reg[28][11]  (.Q (\values[28] [11] ), .CK (n_121_91), .D (sps__n12));
DFF_X1 \values_reg[28][12]  (.Q (\values[28] [12] ), .CK (n_121_91), .D (sps__n57));
DFF_X1 \values_reg[28][13]  (.Q (\values[28] [13] ), .CK (n_121_91), .D (sps__n39));
DFF_X1 \values_reg[28][14]  (.Q (\values[28] [14] ), .CK (n_121_91), .D (sps__n25));
DFF_X1 \values_reg[28][15]  (.Q (\values[28] [15] ), .CK (n_121_91), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[28]_reg  (.GCK (n_121_91), .CK (clk), .E (n_28), .SE (1'b0 ));
DFF_X1 \values_reg[29][0]  (.Q (\values[29] [0] ), .CK (n_121_90), .D (sps__n5));
DFF_X1 \values_reg[29][1]  (.Q (\values[29] [1] ), .CK (n_121_90), .D (sps__n71));
DFF_X1 \values_reg[29][2]  (.Q (\values[29] [2] ), .CK (n_121_90), .D (spc__n159));
DFF_X1 \values_reg[29][3]  (.Q (\values[29] [3] ), .CK (n_121_90), .D (sps__n78));
DFF_X1 \values_reg[29][4]  (.Q (\values[29] [4] ), .CK (n_121_90), .D (sps__n89));
DFF_X1 \values_reg[29][5]  (.Q (\values[29] [5] ), .CK (n_121_90), .D (spc__n132));
DFF_X1 \values_reg[29][6]  (.Q (\values[29] [6] ), .CK (n_121_90), .D (sps__n118));
DFF_X1 \values_reg[29][7]  (.Q (\values[29] [7] ), .CK (n_121_90), .D (spc__n127));
DFF_X1 \values_reg[29][8]  (.Q (\values[29] [8] ), .CK (n_121_90), .D (sps__n97));
DFF_X1 \values_reg[29][9]  (.Q (\values[29] [9] ), .CK (n_121_90), .D (sps__n109));
DFF_X1 \values_reg[29][10]  (.Q (\values[29] [10] ), .CK (n_121_90), .D (sps__n1));
DFF_X1 \values_reg[29][11]  (.Q (\values[29] [11] ), .CK (n_121_90), .D (sps__n10));
DFF_X1 \values_reg[29][12]  (.Q (\values[29] [12] ), .CK (n_121_90), .D (sps__n52));
DFF_X1 \values_reg[29][13]  (.Q (\values[29] [13] ), .CK (n_121_90), .D (sps__n39));
DFF_X1 \values_reg[29][14]  (.Q (\values[29] [14] ), .CK (n_121_90), .D (sps__n28));
DFF_X1 \values_reg[29][15]  (.Q (\values[29] [15] ), .CK (n_121_90), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[29]_reg  (.GCK (n_121_90), .CK (clk), .E (n_29), .SE (1'b0 ));
DFF_X1 \values_reg[30][0]  (.Q (\values[30] [0] ), .CK (n_121_89), .D (sps__n5));
DFF_X1 \values_reg[30][1]  (.Q (\values[30] [1] ), .CK (n_121_89), .D (sps__n71));
DFF_X1 \values_reg[30][2]  (.Q (\values[30] [2] ), .CK (n_121_89), .D (spc__n159));
DFF_X1 \values_reg[30][3]  (.Q (\values[30] [3] ), .CK (n_121_89), .D (sps__n77));
DFF_X1 \values_reg[30][4]  (.Q (\values[30] [4] ), .CK (n_121_89), .D (sps__n89));
DFF_X1 \values_reg[30][5]  (.Q (\values[30] [5] ), .CK (n_121_89), .D (spc__n132));
DFF_X1 \values_reg[30][6]  (.Q (\values[30] [6] ), .CK (n_121_89), .D (sps__n117));
DFF_X1 \values_reg[30][7]  (.Q (\values[30] [7] ), .CK (n_121_89), .D (spc__n127));
DFF_X1 \values_reg[30][8]  (.Q (\values[30] [8] ), .CK (n_121_89), .D (sps__n97));
DFF_X1 \values_reg[30][9]  (.Q (\values[30] [9] ), .CK (n_121_89), .D (sps__n108));
DFF_X1 \values_reg[30][10]  (.Q (\values[30] [10] ), .CK (n_121_89), .D (sps__n1));
DFF_X1 \values_reg[30][11]  (.Q (\values[30] [11] ), .CK (n_121_89), .D (sps__n11));
DFF_X1 \values_reg[30][12]  (.Q (\values[30] [12] ), .CK (n_121_89), .D (sps__n57));
DFF_X1 \values_reg[30][13]  (.Q (\values[30] [13] ), .CK (n_121_89), .D (sps__n39));
DFF_X1 \values_reg[30][14]  (.Q (\values[30] [14] ), .CK (n_121_89), .D (sps__n25));
DFF_X1 \values_reg[30][15]  (.Q (\values[30] [15] ), .CK (n_121_89), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[30]_reg  (.GCK (n_121_89), .CK (clk), .E (n_30), .SE (1'b0 ));
DFF_X1 \values_reg[31][0]  (.Q (\values[31] [0] ), .CK (n_121_88), .D (sps__n5));
DFF_X1 \values_reg[31][1]  (.Q (\values[31] [1] ), .CK (n_121_88), .D (sps__n71));
DFF_X1 \values_reg[31][2]  (.Q (\values[31] [2] ), .CK (n_121_88), .D (spc__n157));
DFF_X1 \values_reg[31][3]  (.Q (\values[31] [3] ), .CK (n_121_88), .D (sps__n78));
DFF_X1 \values_reg[31][4]  (.Q (\values[31] [4] ), .CK (n_121_88), .D (sps__n89));
DFF_X1 \values_reg[31][5]  (.Q (\values[31] [5] ), .CK (n_121_88), .D (spc__n132));
DFF_X1 \values_reg[31][6]  (.Q (\values[31] [6] ), .CK (n_121_88), .D (sps__n118));
DFF_X1 \values_reg[31][7]  (.Q (\values[31] [7] ), .CK (n_121_88), .D (spc__n127));
DFF_X1 \values_reg[31][8]  (.Q (\values[31] [8] ), .CK (n_121_88), .D (sps__n97));
DFF_X1 \values_reg[31][9]  (.Q (\values[31] [9] ), .CK (n_121_88), .D (sps__n109));
DFF_X1 \values_reg[31][10]  (.Q (\values[31] [10] ), .CK (n_121_88), .D (sps__n1));
DFF_X1 \values_reg[31][11]  (.Q (\values[31] [11] ), .CK (n_121_88), .D (sps__n10));
DFF_X1 \values_reg[31][12]  (.Q (\values[31] [12] ), .CK (n_121_88), .D (sps__n52));
DFF_X1 \values_reg[31][13]  (.Q (\values[31] [13] ), .CK (n_121_88), .D (sps__n37));
DFF_X1 \values_reg[31][14]  (.Q (\values[31] [14] ), .CK (n_121_88), .D (sps__n28));
DFF_X1 \values_reg[31][15]  (.Q (\values[31] [15] ), .CK (n_121_88), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[31]_reg  (.GCK (n_121_88), .CK (clk), .E (n_31), .SE (1'b0 ));
DFF_X1 \values_reg[32][0]  (.Q (\values[32] [0] ), .CK (n_121_87), .D (sps__n5));
DFF_X1 \values_reg[32][1]  (.Q (\values[32] [1] ), .CK (n_121_87), .D (sps__n71));
DFF_X1 \values_reg[32][2]  (.Q (\values[32] [2] ), .CK (n_121_87), .D (spc__n157));
DFF_X1 \values_reg[32][3]  (.Q (\values[32] [3] ), .CK (n_121_87), .D (sps__n79));
DFF_X1 \values_reg[32][4]  (.Q (\values[32] [4] ), .CK (n_121_87), .D (sps__n89));
DFF_X1 \values_reg[32][5]  (.Q (\values[32] [5] ), .CK (n_121_87), .D (spc__n132));
DFF_X1 \values_reg[32][6]  (.Q (\values[32] [6] ), .CK (n_121_87), .D (sps__n118));
DFF_X1 \values_reg[32][7]  (.Q (\values[32] [7] ), .CK (n_121_87), .D (spc__n126));
DFF_X1 \values_reg[32][8]  (.Q (\values[32] [8] ), .CK (n_121_87), .D (sps__n97));
DFF_X1 \values_reg[32][9]  (.Q (\values[32] [9] ), .CK (n_121_87), .D (sps__n110));
DFF_X1 \values_reg[32][10]  (.Q (\values[32] [10] ), .CK (n_121_87), .D (sps__n1));
DFF_X1 \values_reg[32][11]  (.Q (\values[32] [11] ), .CK (n_121_87), .D (sps__n14));
DFF_X1 \values_reg[32][12]  (.Q (\values[32] [12] ), .CK (n_121_87), .D (sps__n55));
DFF_X1 \values_reg[32][13]  (.Q (\values[32] [13] ), .CK (n_121_87), .D (sps__n38));
DFF_X1 \values_reg[32][14]  (.Q (\values[32] [14] ), .CK (n_121_87), .D (sps__n28));
DFF_X1 \values_reg[32][15]  (.Q (\values[32] [15] ), .CK (n_121_87), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[32]_reg  (.GCK (n_121_87), .CK (clk), .E (n_32), .SE (1'b0 ));
DFF_X1 \values_reg[33][0]  (.Q (\values[33] [0] ), .CK (n_121_86), .D (sps__n5));
DFF_X1 \values_reg[33][1]  (.Q (\values[33] [1] ), .CK (n_121_86), .D (sps__n71));
DFF_X1 \values_reg[33][2]  (.Q (\values[33] [2] ), .CK (n_121_86), .D (spc__n158));
DFF_X1 \values_reg[33][3]  (.Q (\values[33] [3] ), .CK (n_121_86), .D (sps__n79));
DFF_X1 \values_reg[33][4]  (.Q (\values[33] [4] ), .CK (n_121_86), .D (sps__n89));
DFF_X1 \values_reg[33][5]  (.Q (\values[33] [5] ), .CK (n_121_86), .D (spc__n132));
DFF_X1 \values_reg[33][6]  (.Q (\values[33] [6] ), .CK (n_121_86), .D (sps__n119));
DFF_X1 \values_reg[33][7]  (.Q (\values[33] [7] ), .CK (n_121_86), .D (spc__n126));
DFF_X1 \values_reg[33][8]  (.Q (\values[33] [8] ), .CK (n_121_86), .D (sps__n97));
DFF_X1 \values_reg[33][9]  (.Q (\values[33] [9] ), .CK (n_121_86), .D (sps__n110));
DFF_X1 \values_reg[33][10]  (.Q (\values[33] [10] ), .CK (n_121_86), .D (sps__n1));
DFF_X1 \values_reg[33][11]  (.Q (\values[33] [11] ), .CK (n_121_86), .D (sps__n14));
DFF_X1 \values_reg[33][12]  (.Q (\values[33] [12] ), .CK (n_121_86), .D (sps__n55));
DFF_X1 \values_reg[33][13]  (.Q (\values[33] [13] ), .CK (n_121_86), .D (sps__n38));
DFF_X1 \values_reg[33][14]  (.Q (\values[33] [14] ), .CK (n_121_86), .D (sps__n28));
DFF_X1 \values_reg[33][15]  (.Q (\values[33] [15] ), .CK (n_121_86), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[33]_reg  (.GCK (n_121_86), .CK (clk), .E (n_33), .SE (1'b0 ));
DFF_X1 \values_reg[34][0]  (.Q (\values[34] [0] ), .CK (n_121_85), .D (sps__n5));
DFF_X1 \values_reg[34][1]  (.Q (\values[34] [1] ), .CK (n_121_85), .D (sps__n71));
DFF_X1 \values_reg[34][2]  (.Q (\values[34] [2] ), .CK (n_121_85), .D (spc__n158));
DFF_X1 \values_reg[34][3]  (.Q (\values[34] [3] ), .CK (n_121_85), .D (sps__n79));
DFF_X1 \values_reg[34][4]  (.Q (\values[34] [4] ), .CK (n_121_85), .D (sps__n89));
DFF_X1 \values_reg[34][5]  (.Q (\values[34] [5] ), .CK (n_121_85), .D (spc__n132));
DFF_X1 \values_reg[34][6]  (.Q (\values[34] [6] ), .CK (n_121_85), .D (sps__n119));
DFF_X1 \values_reg[34][7]  (.Q (\values[34] [7] ), .CK (n_121_85), .D (spc__n126));
DFF_X1 \values_reg[34][8]  (.Q (\values[34] [8] ), .CK (n_121_85), .D (sps__n97));
DFF_X1 \values_reg[34][9]  (.Q (\values[34] [9] ), .CK (n_121_85), .D (sps__n110));
DFF_X1 \values_reg[34][10]  (.Q (\values[34] [10] ), .CK (n_121_85), .D (sps__n1));
DFF_X1 \values_reg[34][11]  (.Q (\values[34] [11] ), .CK (n_121_85), .D (sps__n14));
DFF_X1 \values_reg[34][12]  (.Q (\values[34] [12] ), .CK (n_121_85), .D (sps__n55));
DFF_X1 \values_reg[34][13]  (.Q (\values[34] [13] ), .CK (n_121_85), .D (sps__n38));
DFF_X1 \values_reg[34][14]  (.Q (\values[34] [14] ), .CK (n_121_85), .D (sps__n28));
DFF_X1 \values_reg[34][15]  (.Q (\values[34] [15] ), .CK (n_121_85), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[34]_reg  (.GCK (n_121_85), .CK (clk), .E (n_34), .SE (1'b0 ));
DFF_X1 \values_reg[35][0]  (.Q (\values[35] [0] ), .CK (n_121_84), .D (sps__n5));
DFF_X1 \values_reg[35][1]  (.Q (\values[35] [1] ), .CK (n_121_84), .D (sps__n71));
DFF_X1 \values_reg[35][2]  (.Q (\values[35] [2] ), .CK (n_121_84), .D (spc__n158));
DFF_X1 \values_reg[35][3]  (.Q (\values[35] [3] ), .CK (n_121_84), .D (sps__n79));
DFF_X1 \values_reg[35][4]  (.Q (\values[35] [4] ), .CK (n_121_84), .D (sps__n89));
DFF_X1 \values_reg[35][5]  (.Q (\values[35] [5] ), .CK (n_121_84), .D (spc__n132));
DFF_X1 \values_reg[35][6]  (.Q (\values[35] [6] ), .CK (n_121_84), .D (sps__n119));
DFF_X1 \values_reg[35][7]  (.Q (\values[35] [7] ), .CK (n_121_84), .D (spc__n127));
DFF_X1 \values_reg[35][8]  (.Q (\values[35] [8] ), .CK (n_121_84), .D (sps__n97));
DFF_X1 \values_reg[35][9]  (.Q (\values[35] [9] ), .CK (n_121_84), .D (sps__n108));
DFF_X1 \values_reg[35][10]  (.Q (\values[35] [10] ), .CK (n_121_84), .D (sps__n1));
DFF_X1 \values_reg[35][11]  (.Q (\values[35] [11] ), .CK (n_121_84), .D (sps__n11));
DFF_X1 \values_reg[35][12]  (.Q (\values[35] [12] ), .CK (n_121_84), .D (sps__n57));
DFF_X1 \values_reg[35][13]  (.Q (\values[35] [13] ), .CK (n_121_84), .D (sps__n38));
DFF_X1 \values_reg[35][14]  (.Q (\values[35] [14] ), .CK (n_121_84), .D (sps__n28));
DFF_X1 \values_reg[35][15]  (.Q (\values[35] [15] ), .CK (n_121_84), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[35]_reg  (.GCK (n_121_84), .CK (clk), .E (n_35), .SE (1'b0 ));
DFF_X1 \values_reg[36][0]  (.Q (\values[36] [0] ), .CK (n_121_83), .D (sps__n5));
DFF_X1 \values_reg[36][1]  (.Q (\values[36] [1] ), .CK (n_121_83), .D (sps__n71));
DFF_X1 \values_reg[36][2]  (.Q (\values[36] [2] ), .CK (n_121_83), .D (spc__n158));
DFF_X1 \values_reg[36][3]  (.Q (\values[36] [3] ), .CK (n_121_83), .D (sps__n79));
DFF_X1 \values_reg[36][4]  (.Q (\values[36] [4] ), .CK (n_121_83), .D (sps__n89));
DFF_X1 \values_reg[36][5]  (.Q (\values[36] [5] ), .CK (n_121_83), .D (spc__n132));
DFF_X1 \values_reg[36][6]  (.Q (\values[36] [6] ), .CK (n_121_83), .D (sps__n119));
DFF_X1 \values_reg[36][7]  (.Q (\values[36] [7] ), .CK (n_121_83), .D (spc__n126));
DFF_X1 \values_reg[36][8]  (.Q (\values[36] [8] ), .CK (n_121_83), .D (sps__n97));
DFF_X1 \values_reg[36][9]  (.Q (\values[36] [9] ), .CK (n_121_83), .D (sps__n110));
DFF_X1 \values_reg[36][10]  (.Q (\values[36] [10] ), .CK (n_121_83), .D (sps__n1));
DFF_X1 \values_reg[36][11]  (.Q (\values[36] [11] ), .CK (n_121_83), .D (sps__n14));
DFF_X1 \values_reg[36][12]  (.Q (\values[36] [12] ), .CK (n_121_83), .D (sps__n55));
DFF_X1 \values_reg[36][13]  (.Q (\values[36] [13] ), .CK (n_121_83), .D (sps__n38));
DFF_X1 \values_reg[36][14]  (.Q (\values[36] [14] ), .CK (n_121_83), .D (sps__n28));
DFF_X1 \values_reg[36][15]  (.Q (\values[36] [15] ), .CK (n_121_83), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[36]_reg  (.GCK (n_121_83), .CK (clk), .E (n_36), .SE (1'b0 ));
DFF_X1 \values_reg[37][0]  (.Q (\values[37] [0] ), .CK (n_121_82), .D (sps__n5));
DFF_X1 \values_reg[37][1]  (.Q (\values[37] [1] ), .CK (n_121_82), .D (sps__n71));
DFF_X1 \values_reg[37][2]  (.Q (\values[37] [2] ), .CK (n_121_82), .D (spc__n158));
DFF_X1 \values_reg[37][3]  (.Q (\values[37] [3] ), .CK (n_121_82), .D (sps__n79));
DFF_X1 \values_reg[37][4]  (.Q (\values[37] [4] ), .CK (n_121_82), .D (sps__n89));
DFF_X1 \values_reg[37][5]  (.Q (\values[37] [5] ), .CK (n_121_82), .D (spc__n132));
DFF_X1 \values_reg[37][6]  (.Q (\values[37] [6] ), .CK (n_121_82), .D (sps__n119));
DFF_X1 \values_reg[37][7]  (.Q (\values[37] [7] ), .CK (n_121_82), .D (spc__n126));
DFF_X1 \values_reg[37][8]  (.Q (\values[37] [8] ), .CK (n_121_82), .D (sps__n97));
DFF_X1 \values_reg[37][9]  (.Q (\values[37] [9] ), .CK (n_121_82), .D (sps__n110));
DFF_X1 \values_reg[37][10]  (.Q (\values[37] [10] ), .CK (n_121_82), .D (sps__n1));
DFF_X1 \values_reg[37][11]  (.Q (\values[37] [11] ), .CK (n_121_82), .D (sps__n14));
DFF_X1 \values_reg[37][12]  (.Q (\values[37] [12] ), .CK (n_121_82), .D (sps__n55));
DFF_X1 \values_reg[37][13]  (.Q (\values[37] [13] ), .CK (n_121_82), .D (sps__n38));
DFF_X1 \values_reg[37][14]  (.Q (\values[37] [14] ), .CK (n_121_82), .D (sps__n28));
DFF_X1 \values_reg[37][15]  (.Q (\values[37] [15] ), .CK (n_121_82), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[37]_reg  (.GCK (n_121_82), .CK (clk), .E (n_37), .SE (1'b0 ));
DFF_X1 \values_reg[38][0]  (.Q (\values[38] [0] ), .CK (n_121_81), .D (sps__n5));
DFF_X1 \values_reg[38][1]  (.Q (\values[38] [1] ), .CK (n_121_81), .D (sps__n71));
DFF_X1 \values_reg[38][2]  (.Q (\values[38] [2] ), .CK (n_121_81), .D (spc__n158));
DFF_X1 \values_reg[38][3]  (.Q (\values[38] [3] ), .CK (n_121_81), .D (sps__n79));
DFF_X1 \values_reg[38][4]  (.Q (\values[38] [4] ), .CK (n_121_81), .D (sps__n89));
DFF_X1 \values_reg[38][5]  (.Q (\values[38] [5] ), .CK (n_121_81), .D (spc__n132));
DFF_X1 \values_reg[38][6]  (.Q (\values[38] [6] ), .CK (n_121_81), .D (sps__n119));
DFF_X1 \values_reg[38][7]  (.Q (\values[38] [7] ), .CK (n_121_81), .D (spc__n126));
DFF_X1 \values_reg[38][8]  (.Q (\values[38] [8] ), .CK (n_121_81), .D (sps__n97));
DFF_X1 \values_reg[38][9]  (.Q (\values[38] [9] ), .CK (n_121_81), .D (sps__n108));
DFF_X1 \values_reg[38][10]  (.Q (\values[38] [10] ), .CK (n_121_81), .D (sps__n1));
DFF_X1 \values_reg[38][11]  (.Q (\values[38] [11] ), .CK (n_121_81), .D (sps__n14));
DFF_X1 \values_reg[38][12]  (.Q (\values[38] [12] ), .CK (n_121_81), .D (sps__n55));
DFF_X1 \values_reg[38][13]  (.Q (\values[38] [13] ), .CK (n_121_81), .D (sps__n38));
DFF_X1 \values_reg[38][14]  (.Q (\values[38] [14] ), .CK (n_121_81), .D (sps__n28));
DFF_X1 \values_reg[38][15]  (.Q (\values[38] [15] ), .CK (n_121_81), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[38]_reg  (.GCK (n_121_81), .CK (clk), .E (n_38), .SE (1'b0 ));
DFF_X1 \values_reg[39][0]  (.Q (\values[39] [0] ), .CK (n_121_80), .D (sps__n5));
DFF_X1 \values_reg[39][1]  (.Q (\values[39] [1] ), .CK (n_121_80), .D (sps__n71));
DFF_X1 \values_reg[39][2]  (.Q (\values[39] [2] ), .CK (n_121_80), .D (spc__n159));
DFF_X1 \values_reg[39][3]  (.Q (\values[39] [3] ), .CK (n_121_80), .D (sps__n79));
DFF_X1 \values_reg[39][4]  (.Q (\values[39] [4] ), .CK (n_121_80), .D (sps__n89));
DFF_X1 \values_reg[39][5]  (.Q (\values[39] [5] ), .CK (n_121_80), .D (spc__n132));
DFF_X1 \values_reg[39][6]  (.Q (\values[39] [6] ), .CK (n_121_80), .D (sps__n119));
DFF_X1 \values_reg[39][7]  (.Q (\values[39] [7] ), .CK (n_121_80), .D (spc__n127));
DFF_X1 \values_reg[39][8]  (.Q (\values[39] [8] ), .CK (n_121_80), .D (sps__n97));
DFF_X1 \values_reg[39][9]  (.Q (\values[39] [9] ), .CK (n_121_80), .D (sps__n108));
DFF_X1 \values_reg[39][10]  (.Q (\values[39] [10] ), .CK (n_121_80), .D (sps__n1));
DFF_X1 \values_reg[39][11]  (.Q (\values[39] [11] ), .CK (n_121_80), .D (sps__n11));
DFF_X1 \values_reg[39][12]  (.Q (\values[39] [12] ), .CK (n_121_80), .D (sps__n55));
DFF_X1 \values_reg[39][13]  (.Q (\values[39] [13] ), .CK (n_121_80), .D (sps__n38));
DFF_X1 \values_reg[39][14]  (.Q (\values[39] [14] ), .CK (n_121_80), .D (sps__n28));
DFF_X1 \values_reg[39][15]  (.Q (\values[39] [15] ), .CK (n_121_80), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[39]_reg  (.GCK (n_121_80), .CK (clk), .E (n_39), .SE (1'b0 ));
DFF_X1 \values_reg[40][0]  (.Q (\values[40] [0] ), .CK (n_121_79), .D (sps__n5));
DFF_X1 \values_reg[40][1]  (.Q (\values[40] [1] ), .CK (n_121_79), .D (sps__n71));
DFF_X1 \values_reg[40][2]  (.Q (\values[40] [2] ), .CK (n_121_79), .D (spc__n158));
DFF_X1 \values_reg[40][3]  (.Q (\values[40] [3] ), .CK (n_121_79), .D (sps__n79));
DFF_X1 \values_reg[40][4]  (.Q (\values[40] [4] ), .CK (n_121_79), .D (sps__n89));
DFF_X1 \values_reg[40][5]  (.Q (\values[40] [5] ), .CK (n_121_79), .D (spc__n132));
DFF_X1 \values_reg[40][6]  (.Q (\values[40] [6] ), .CK (n_121_79), .D (sps__n118));
DFF_X1 \values_reg[40][7]  (.Q (\values[40] [7] ), .CK (n_121_79), .D (spc__n126));
DFF_X1 \values_reg[40][8]  (.Q (\values[40] [8] ), .CK (n_121_79), .D (sps__n97));
DFF_X1 \values_reg[40][9]  (.Q (\values[40] [9] ), .CK (n_121_79), .D (sps__n110));
DFF_X1 \values_reg[40][10]  (.Q (\values[40] [10] ), .CK (n_121_79), .D (sps__n1));
DFF_X1 \values_reg[40][11]  (.Q (\values[40] [11] ), .CK (n_121_79), .D (sps__n14));
DFF_X1 \values_reg[40][12]  (.Q (\values[40] [12] ), .CK (n_121_79), .D (sps__n55));
DFF_X1 \values_reg[40][13]  (.Q (\values[40] [13] ), .CK (n_121_79), .D (sps__n40));
DFF_X1 \values_reg[40][14]  (.Q (\values[40] [14] ), .CK (n_121_79), .D (sps__n28));
DFF_X1 \values_reg[40][15]  (.Q (\values[40] [15] ), .CK (n_121_79), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[40]_reg  (.GCK (n_121_79), .CK (clk), .E (n_40), .SE (1'b0 ));
DFF_X1 \values_reg[41][0]  (.Q (\values[41] [0] ), .CK (n_121_78), .D (sps__n5));
DFF_X1 \values_reg[41][1]  (.Q (\values[41] [1] ), .CK (n_121_78), .D (sps__n71));
DFF_X1 \values_reg[41][2]  (.Q (\values[41] [2] ), .CK (n_121_78), .D (spc__n157));
DFF_X1 \values_reg[41][3]  (.Q (\values[41] [3] ), .CK (n_121_78), .D (sps__n79));
DFF_X1 \values_reg[41][4]  (.Q (\values[41] [4] ), .CK (n_121_78), .D (sps__n89));
DFF_X1 \values_reg[41][5]  (.Q (\values[41] [5] ), .CK (n_121_78), .D (spc__n132));
DFF_X1 \values_reg[41][6]  (.Q (\values[41] [6] ), .CK (n_121_78), .D (sps__n118));
DFF_X1 \values_reg[41][7]  (.Q (\values[41] [7] ), .CK (n_121_78), .D (spc__n126));
DFF_X1 \values_reg[41][8]  (.Q (\values[41] [8] ), .CK (n_121_78), .D (sps__n97));
DFF_X1 \values_reg[41][9]  (.Q (\values[41] [9] ), .CK (n_121_78), .D (sps__n110));
DFF_X1 \values_reg[41][10]  (.Q (\values[41] [10] ), .CK (n_121_78), .D (sps__n1));
DFF_X1 \values_reg[41][11]  (.Q (\values[41] [11] ), .CK (n_121_78), .D (sps__n14));
DFF_X1 \values_reg[41][12]  (.Q (\values[41] [12] ), .CK (n_121_78), .D (sps__n55));
DFF_X1 \values_reg[41][13]  (.Q (\values[41] [13] ), .CK (n_121_78), .D (sps__n40));
DFF_X1 \values_reg[41][14]  (.Q (\values[41] [14] ), .CK (n_121_78), .D (sps__n28));
DFF_X1 \values_reg[41][15]  (.Q (\values[41] [15] ), .CK (n_121_78), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[41]_reg  (.GCK (n_121_78), .CK (clk), .E (n_41), .SE (1'b0 ));
DFF_X1 \values_reg[42][0]  (.Q (\values[42] [0] ), .CK (n_121_77), .D (sps__n5));
DFF_X1 \values_reg[42][1]  (.Q (\values[42] [1] ), .CK (n_121_77), .D (sps__n71));
DFF_X1 \values_reg[42][2]  (.Q (\values[42] [2] ), .CK (n_121_77), .D (spc__n158));
DFF_X1 \values_reg[42][3]  (.Q (\values[42] [3] ), .CK (n_121_77), .D (sps__n79));
DFF_X1 \values_reg[42][4]  (.Q (\values[42] [4] ), .CK (n_121_77), .D (sps__n89));
DFF_X1 \values_reg[42][5]  (.Q (\values[42] [5] ), .CK (n_121_77), .D (spc__n132));
DFF_X1 \values_reg[42][6]  (.Q (\values[42] [6] ), .CK (n_121_77), .D (sps__n119));
DFF_X1 \values_reg[42][7]  (.Q (\values[42] [7] ), .CK (n_121_77), .D (spc__n126));
DFF_X1 \values_reg[42][8]  (.Q (\values[42] [8] ), .CK (n_121_77), .D (sps__n97));
DFF_X1 \values_reg[42][9]  (.Q (\values[42] [9] ), .CK (n_121_77), .D (sps__n110));
DFF_X1 \values_reg[42][10]  (.Q (\values[42] [10] ), .CK (n_121_77), .D (sps__n1));
DFF_X1 \values_reg[42][11]  (.Q (\values[42] [11] ), .CK (n_121_77), .D (sps__n14));
DFF_X1 \values_reg[42][12]  (.Q (\values[42] [12] ), .CK (n_121_77), .D (sps__n55));
DFF_X1 \values_reg[42][13]  (.Q (\values[42] [13] ), .CK (n_121_77), .D (sps__n40));
DFF_X1 \values_reg[42][14]  (.Q (\values[42] [14] ), .CK (n_121_77), .D (sps__n28));
DFF_X1 \values_reg[42][15]  (.Q (\values[42] [15] ), .CK (n_121_77), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[42]_reg  (.GCK (n_121_77), .CK (clk), .E (n_42), .SE (1'b0 ));
DFF_X1 \values_reg[43][0]  (.Q (\values[43] [0] ), .CK (n_121_76), .D (sps__n5));
DFF_X1 \values_reg[43][1]  (.Q (\values[43] [1] ), .CK (n_121_76), .D (sps__n71));
DFF_X1 \values_reg[43][2]  (.Q (\values[43] [2] ), .CK (n_121_76), .D (spc__n157));
DFF_X1 \values_reg[43][3]  (.Q (\values[43] [3] ), .CK (n_121_76), .D (sps__n79));
DFF_X1 \values_reg[43][4]  (.Q (\values[43] [4] ), .CK (n_121_76), .D (sps__n89));
DFF_X1 \values_reg[43][5]  (.Q (\values[43] [5] ), .CK (n_121_76), .D (spc__n132));
DFF_X1 \values_reg[43][6]  (.Q (\values[43] [6] ), .CK (n_121_76), .D (sps__n119));
DFF_X1 \values_reg[43][7]  (.Q (\values[43] [7] ), .CK (n_121_76), .D (spc__n126));
DFF_X1 \values_reg[43][8]  (.Q (\values[43] [8] ), .CK (n_121_76), .D (sps__n97));
DFF_X1 \values_reg[43][9]  (.Q (\values[43] [9] ), .CK (n_121_76), .D (sps__n109));
DFF_X1 \values_reg[43][10]  (.Q (\values[43] [10] ), .CK (n_121_76), .D (sps__n1));
DFF_X1 \values_reg[43][11]  (.Q (\values[43] [11] ), .CK (n_121_76), .D (sps__n14));
DFF_X1 \values_reg[43][12]  (.Q (\values[43] [12] ), .CK (n_121_76), .D (sps__n55));
DFF_X1 \values_reg[43][13]  (.Q (\values[43] [13] ), .CK (n_121_76), .D (sps__n40));
DFF_X1 \values_reg[43][14]  (.Q (\values[43] [14] ), .CK (n_121_76), .D (sps__n28));
DFF_X1 \values_reg[43][15]  (.Q (\values[43] [15] ), .CK (n_121_76), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[43]_reg  (.GCK (n_121_76), .CK (clk), .E (n_43), .SE (1'b0 ));
DFF_X1 \values_reg[44][0]  (.Q (\values[44] [0] ), .CK (n_121_75), .D (sps__n5));
DFF_X1 \values_reg[44][1]  (.Q (\values[44] [1] ), .CK (n_121_75), .D (sps__n71));
DFF_X1 \values_reg[44][2]  (.Q (\values[44] [2] ), .CK (n_121_75), .D (spc__n157));
DFF_X1 \values_reg[44][3]  (.Q (\values[44] [3] ), .CK (n_121_75), .D (sps__n79));
DFF_X1 \values_reg[44][4]  (.Q (\values[44] [4] ), .CK (n_121_75), .D (sps__n89));
DFF_X1 \values_reg[44][5]  (.Q (\values[44] [5] ), .CK (n_121_75), .D (spc__n132));
DFF_X1 \values_reg[44][6]  (.Q (\values[44] [6] ), .CK (n_121_75), .D (sps__n118));
DFF_X1 \values_reg[44][7]  (.Q (\values[44] [7] ), .CK (n_121_75), .D (spc__n126));
DFF_X1 \values_reg[44][8]  (.Q (\values[44] [8] ), .CK (n_121_75), .D (sps__n97));
DFF_X1 \values_reg[44][9]  (.Q (\values[44] [9] ), .CK (n_121_75), .D (sps__n109));
DFF_X1 \values_reg[44][10]  (.Q (\values[44] [10] ), .CK (n_121_75), .D (sps__n1));
DFF_X1 \values_reg[44][11]  (.Q (\values[44] [11] ), .CK (n_121_75), .D (sps__n14));
DFF_X1 \values_reg[44][12]  (.Q (\values[44] [12] ), .CK (n_121_75), .D (sps__n55));
DFF_X1 \values_reg[44][13]  (.Q (\values[44] [13] ), .CK (n_121_75), .D (sps__n40));
DFF_X1 \values_reg[44][14]  (.Q (\values[44] [14] ), .CK (n_121_75), .D (sps__n28));
DFF_X1 \values_reg[44][15]  (.Q (\values[44] [15] ), .CK (n_121_75), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[44]_reg  (.GCK (n_121_75), .CK (clk), .E (n_44), .SE (1'b0 ));
DFF_X1 \values_reg[45][0]  (.Q (\values[45] [0] ), .CK (n_121_74), .D (sps__n5));
DFF_X1 \values_reg[45][1]  (.Q (\values[45] [1] ), .CK (n_121_74), .D (sps__n71));
DFF_X1 \values_reg[45][2]  (.Q (\values[45] [2] ), .CK (n_121_74), .D (spc__n157));
DFF_X1 \values_reg[45][3]  (.Q (\values[45] [3] ), .CK (n_121_74), .D (sps__n79));
DFF_X1 \values_reg[45][4]  (.Q (\values[45] [4] ), .CK (n_121_74), .D (sps__n89));
DFF_X1 \values_reg[45][5]  (.Q (\values[45] [5] ), .CK (n_121_74), .D (spc__n132));
DFF_X1 \values_reg[45][6]  (.Q (\values[45] [6] ), .CK (n_121_74), .D (sps__n118));
DFF_X1 \values_reg[45][7]  (.Q (\values[45] [7] ), .CK (n_121_74), .D (spc__n126));
DFF_X1 \values_reg[45][8]  (.Q (\values[45] [8] ), .CK (n_121_74), .D (sps__n97));
DFF_X1 \values_reg[45][9]  (.Q (\values[45] [9] ), .CK (n_121_74), .D (sps__n109));
DFF_X1 \values_reg[45][10]  (.Q (\values[45] [10] ), .CK (n_121_74), .D (sps__n1));
DFF_X1 \values_reg[45][11]  (.Q (\values[45] [11] ), .CK (n_121_74), .D (sps__n14));
DFF_X1 \values_reg[45][12]  (.Q (\values[45] [12] ), .CK (n_121_74), .D (sps__n55));
DFF_X1 \values_reg[45][13]  (.Q (\values[45] [13] ), .CK (n_121_74), .D (sps__n40));
DFF_X1 \values_reg[45][14]  (.Q (\values[45] [14] ), .CK (n_121_74), .D (sps__n28));
DFF_X1 \values_reg[45][15]  (.Q (\values[45] [15] ), .CK (n_121_74), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[45]_reg  (.GCK (n_121_74), .CK (clk), .E (n_45), .SE (1'b0 ));
DFF_X1 \values_reg[46][0]  (.Q (\values[46] [0] ), .CK (n_121_73), .D (sps__n5));
DFF_X1 \values_reg[46][1]  (.Q (\values[46] [1] ), .CK (n_121_73), .D (sps__n71));
DFF_X1 \values_reg[46][2]  (.Q (\values[46] [2] ), .CK (n_121_73), .D (spc__n157));
DFF_X1 \values_reg[46][3]  (.Q (\values[46] [3] ), .CK (n_121_73), .D (sps__n79));
DFF_X1 \values_reg[46][4]  (.Q (\values[46] [4] ), .CK (n_121_73), .D (sps__n89));
DFF_X1 \values_reg[46][5]  (.Q (\values[46] [5] ), .CK (n_121_73), .D (spc__n132));
DFF_X1 \values_reg[46][6]  (.Q (\values[46] [6] ), .CK (n_121_73), .D (sps__n118));
DFF_X1 \values_reg[46][7]  (.Q (\values[46] [7] ), .CK (n_121_73), .D (spc__n126));
DFF_X1 \values_reg[46][8]  (.Q (\values[46] [8] ), .CK (n_121_73), .D (sps__n97));
DFF_X1 \values_reg[46][9]  (.Q (\values[46] [9] ), .CK (n_121_73), .D (sps__n109));
DFF_X1 \values_reg[46][10]  (.Q (\values[46] [10] ), .CK (n_121_73), .D (sps__n1));
DFF_X1 \values_reg[46][11]  (.Q (\values[46] [11] ), .CK (n_121_73), .D (sps__n14));
DFF_X1 \values_reg[46][12]  (.Q (\values[46] [12] ), .CK (n_121_73), .D (sps__n55));
DFF_X1 \values_reg[46][13]  (.Q (\values[46] [13] ), .CK (n_121_73), .D (sps__n40));
DFF_X1 \values_reg[46][14]  (.Q (\values[46] [14] ), .CK (n_121_73), .D (sps__n28));
DFF_X1 \values_reg[46][15]  (.Q (\values[46] [15] ), .CK (n_121_73), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[46]_reg  (.GCK (n_121_73), .CK (clk), .E (n_46), .SE (1'b0 ));
DFF_X1 \values_reg[47][0]  (.Q (\values[47] [0] ), .CK (n_121_72), .D (sps__n5));
DFF_X1 \values_reg[47][1]  (.Q (\values[47] [1] ), .CK (n_121_72), .D (sps__n71));
DFF_X1 \values_reg[47][2]  (.Q (\values[47] [2] ), .CK (n_121_72), .D (spc__n157));
DFF_X1 \values_reg[47][3]  (.Q (\values[47] [3] ), .CK (n_121_72), .D (sps__n79));
DFF_X1 \values_reg[47][4]  (.Q (\values[47] [4] ), .CK (n_121_72), .D (sps__n89));
DFF_X1 \values_reg[47][5]  (.Q (\values[47] [5] ), .CK (n_121_72), .D (spc__n132));
DFF_X1 \values_reg[47][6]  (.Q (\values[47] [6] ), .CK (n_121_72), .D (sps__n119));
DFF_X1 \values_reg[47][7]  (.Q (\values[47] [7] ), .CK (n_121_72), .D (spc__n126));
DFF_X1 \values_reg[47][8]  (.Q (\values[47] [8] ), .CK (n_121_72), .D (sps__n97));
DFF_X1 \values_reg[47][9]  (.Q (\values[47] [9] ), .CK (n_121_72), .D (sps__n109));
DFF_X1 \values_reg[47][10]  (.Q (\values[47] [10] ), .CK (n_121_72), .D (sps__n1));
DFF_X1 \values_reg[47][11]  (.Q (\values[47] [11] ), .CK (n_121_72), .D (sps__n14));
DFF_X1 \values_reg[47][12]  (.Q (\values[47] [12] ), .CK (n_121_72), .D (sps__n55));
DFF_X1 \values_reg[47][13]  (.Q (\values[47] [13] ), .CK (n_121_72), .D (sps__n40));
DFF_X1 \values_reg[47][14]  (.Q (\values[47] [14] ), .CK (n_121_72), .D (sps__n28));
DFF_X1 \values_reg[47][15]  (.Q (\values[47] [15] ), .CK (n_121_72), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[47]_reg  (.GCK (n_121_72), .CK (clk), .E (n_47), .SE (1'b0 ));
DFF_X1 \values_reg[48][0]  (.Q (\values[48] [0] ), .CK (n_121_71), .D (sps__n5));
DFF_X1 \values_reg[48][1]  (.Q (\values[48] [1] ), .CK (n_121_71), .D (sps__n71));
DFF_X1 \values_reg[48][2]  (.Q (\values[48] [2] ), .CK (n_121_71), .D (spc__n157));
DFF_X1 \values_reg[48][3]  (.Q (\values[48] [3] ), .CK (n_121_71), .D (sps__n79));
DFF_X1 \values_reg[48][4]  (.Q (\values[48] [4] ), .CK (n_121_71), .D (sps__n89));
DFF_X1 \values_reg[48][5]  (.Q (\values[48] [5] ), .CK (n_121_71), .D (spc__n132));
DFF_X1 \values_reg[48][6]  (.Q (\values[48] [6] ), .CK (n_121_71), .D (sps__n119));
DFF_X1 \values_reg[48][7]  (.Q (\values[48] [7] ), .CK (n_121_71), .D (spc__n126));
DFF_X1 \values_reg[48][8]  (.Q (\values[48] [8] ), .CK (n_121_71), .D (sps__n97));
DFF_X1 \values_reg[48][9]  (.Q (\values[48] [9] ), .CK (n_121_71), .D (sps__n109));
DFF_X1 \values_reg[48][10]  (.Q (\values[48] [10] ), .CK (n_121_71), .D (sps__n1));
DFF_X1 \values_reg[48][11]  (.Q (\values[48] [11] ), .CK (n_121_71), .D (sps__n14));
DFF_X1 \values_reg[48][12]  (.Q (\values[48] [12] ), .CK (n_121_71), .D (sps__n55));
DFF_X1 \values_reg[48][13]  (.Q (\values[48] [13] ), .CK (n_121_71), .D (sps__n40));
DFF_X1 \values_reg[48][14]  (.Q (\values[48] [14] ), .CK (n_121_71), .D (sps__n28));
DFF_X1 \values_reg[48][15]  (.Q (\values[48] [15] ), .CK (n_121_71), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[48]_reg  (.GCK (n_121_71), .CK (clk), .E (n_48), .SE (1'b0 ));
DFF_X1 \values_reg[49][0]  (.Q (\values[49] [0] ), .CK (n_121_70), .D (sps__n5));
DFF_X1 \values_reg[49][1]  (.Q (\values[49] [1] ), .CK (n_121_70), .D (sps__n71));
DFF_X1 \values_reg[49][2]  (.Q (\values[49] [2] ), .CK (n_121_70), .D (spc__n157));
DFF_X1 \values_reg[49][3]  (.Q (\values[49] [3] ), .CK (n_121_70), .D (sps__n76));
DFF_X1 \values_reg[49][4]  (.Q (\values[49] [4] ), .CK (n_121_70), .D (sps__n89));
DFF_X1 \values_reg[49][5]  (.Q (\values[49] [5] ), .CK (n_121_70), .D (spc__n132));
DFF_X1 \values_reg[49][6]  (.Q (\values[49] [6] ), .CK (n_121_70), .D (sps__n118));
DFF_X1 \values_reg[49][7]  (.Q (\values[49] [7] ), .CK (n_121_70), .D (spc__n126));
DFF_X1 \values_reg[49][8]  (.Q (\values[49] [8] ), .CK (n_121_70), .D (sps__n97));
DFF_X1 \values_reg[49][9]  (.Q (\values[49] [9] ), .CK (n_121_70), .D (sps__n110));
DFF_X1 \values_reg[49][10]  (.Q (\values[49] [10] ), .CK (n_121_70), .D (sps__n1));
DFF_X1 \values_reg[49][11]  (.Q (\values[49] [11] ), .CK (n_121_70), .D (sps__n14));
DFF_X1 \values_reg[49][12]  (.Q (\values[49] [12] ), .CK (n_121_70), .D (sps__n55));
DFF_X1 \values_reg[49][13]  (.Q (\values[49] [13] ), .CK (n_121_70), .D (sps__n40));
DFF_X1 \values_reg[49][14]  (.Q (\values[49] [14] ), .CK (n_121_70), .D (sps__n28));
DFF_X1 \values_reg[49][15]  (.Q (\values[49] [15] ), .CK (n_121_70), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[49]_reg  (.GCK (n_121_70), .CK (clk), .E (n_49), .SE (1'b0 ));
DFF_X1 \values_reg[50][0]  (.Q (\values[50] [0] ), .CK (n_121_69), .D (sps__n5));
DFF_X1 \values_reg[50][1]  (.Q (\values[50] [1] ), .CK (n_121_69), .D (sps__n71));
DFF_X1 \values_reg[50][2]  (.Q (\values[50] [2] ), .CK (n_121_69), .D (spc__n159));
DFF_X1 \values_reg[50][3]  (.Q (\values[50] [3] ), .CK (n_121_69), .D (sps__n77));
DFF_X1 \values_reg[50][4]  (.Q (\values[50] [4] ), .CK (n_121_69), .D (sps__n89));
DFF_X1 \values_reg[50][5]  (.Q (\values[50] [5] ), .CK (n_121_69), .D (spc__n132));
DFF_X1 \values_reg[50][6]  (.Q (\values[50] [6] ), .CK (n_121_69), .D (sps__n119));
DFF_X1 \values_reg[50][7]  (.Q (\values[50] [7] ), .CK (n_121_69), .D (spc__n127));
DFF_X1 \values_reg[50][8]  (.Q (\values[50] [8] ), .CK (n_121_69), .D (sps__n97));
DFF_X1 \values_reg[50][9]  (.Q (\values[50] [9] ), .CK (n_121_69), .D (sps__n108));
DFF_X1 \values_reg[50][10]  (.Q (\values[50] [10] ), .CK (n_121_69), .D (sps__n1));
DFF_X1 \values_reg[50][11]  (.Q (\values[50] [11] ), .CK (n_121_69), .D (sps__n11));
DFF_X1 \values_reg[50][12]  (.Q (\values[50] [12] ), .CK (n_121_69), .D (sps__n55));
DFF_X1 \values_reg[50][13]  (.Q (\values[50] [13] ), .CK (n_121_69), .D (sps__n38));
DFF_X1 \values_reg[50][14]  (.Q (\values[50] [14] ), .CK (n_121_69), .D (sps__n28));
DFF_X1 \values_reg[50][15]  (.Q (\values[50] [15] ), .CK (n_121_69), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[50]_reg  (.GCK (n_121_69), .CK (clk), .E (n_50), .SE (1'b0 ));
DFF_X1 \values_reg[51][0]  (.Q (\values[51] [0] ), .CK (n_121_68), .D (sps__n5));
DFF_X1 \values_reg[51][1]  (.Q (\values[51] [1] ), .CK (n_121_68), .D (sps__n71));
DFF_X1 \values_reg[51][2]  (.Q (\values[51] [2] ), .CK (n_121_68), .D (spc__n158));
DFF_X1 \values_reg[51][3]  (.Q (\values[51] [3] ), .CK (n_121_68), .D (sps__n79));
DFF_X1 \values_reg[51][4]  (.Q (\values[51] [4] ), .CK (n_121_68), .D (sps__n89));
DFF_X1 \values_reg[51][5]  (.Q (\values[51] [5] ), .CK (n_121_68), .D (spc__n132));
DFF_X1 \values_reg[51][6]  (.Q (\values[51] [6] ), .CK (n_121_68), .D (sps__n119));
DFF_X1 \values_reg[51][7]  (.Q (\values[51] [7] ), .CK (n_121_68), .D (spc__n126));
DFF_X1 \values_reg[51][8]  (.Q (\values[51] [8] ), .CK (n_121_68), .D (sps__n97));
DFF_X1 \values_reg[51][9]  (.Q (\values[51] [9] ), .CK (n_121_68), .D (sps__n108));
DFF_X1 \values_reg[51][10]  (.Q (\values[51] [10] ), .CK (n_121_68), .D (sps__n1));
DFF_X1 \values_reg[51][11]  (.Q (\values[51] [11] ), .CK (n_121_68), .D (sps__n14));
DFF_X1 \values_reg[51][12]  (.Q (\values[51] [12] ), .CK (n_121_68), .D (sps__n55));
DFF_X1 \values_reg[51][13]  (.Q (\values[51] [13] ), .CK (n_121_68), .D (sps__n38));
DFF_X1 \values_reg[51][14]  (.Q (\values[51] [14] ), .CK (n_121_68), .D (sps__n28));
DFF_X1 \values_reg[51][15]  (.Q (\values[51] [15] ), .CK (n_121_68), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[51]_reg  (.GCK (n_121_68), .CK (clk), .E (n_51), .SE (1'b0 ));
DFF_X1 \values_reg[52][0]  (.Q (\values[52] [0] ), .CK (n_121_67), .D (sps__n5));
DFF_X1 \values_reg[52][1]  (.Q (\values[52] [1] ), .CK (n_121_67), .D (sps__n71));
DFF_X1 \values_reg[52][2]  (.Q (\values[52] [2] ), .CK (n_121_67), .D (spc__n157));
DFF_X1 \values_reg[52][3]  (.Q (\values[52] [3] ), .CK (n_121_67), .D (sps__n79));
DFF_X1 \values_reg[52][4]  (.Q (\values[52] [4] ), .CK (n_121_67), .D (sps__n89));
DFF_X1 \values_reg[52][5]  (.Q (\values[52] [5] ), .CK (n_121_67), .D (spc__n132));
DFF_X1 \values_reg[52][6]  (.Q (\values[52] [6] ), .CK (n_121_67), .D (sps__n118));
DFF_X1 \values_reg[52][7]  (.Q (\values[52] [7] ), .CK (n_121_67), .D (spc__n126));
DFF_X1 \values_reg[52][8]  (.Q (\values[52] [8] ), .CK (n_121_67), .D (sps__n97));
DFF_X1 \values_reg[52][9]  (.Q (\values[52] [9] ), .CK (n_121_67), .D (sps__n110));
DFF_X1 \values_reg[52][10]  (.Q (\values[52] [10] ), .CK (n_121_67), .D (sps__n1));
DFF_X1 \values_reg[52][11]  (.Q (\values[52] [11] ), .CK (n_121_67), .D (sps__n12));
DFF_X1 \values_reg[52][12]  (.Q (\values[52] [12] ), .CK (n_121_67), .D (sps__n55));
DFF_X1 \values_reg[52][13]  (.Q (\values[52] [13] ), .CK (n_121_67), .D (sps__n40));
DFF_X1 \values_reg[52][14]  (.Q (\values[52] [14] ), .CK (n_121_67), .D (sps__n28));
DFF_X1 \values_reg[52][15]  (.Q (\values[52] [15] ), .CK (n_121_67), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[52]_reg  (.GCK (n_121_67), .CK (clk), .E (n_52), .SE (1'b0 ));
DFF_X1 \values_reg[53][0]  (.Q (\values[53] [0] ), .CK (n_121_66), .D (sps__n5));
DFF_X1 \values_reg[53][1]  (.Q (\values[53] [1] ), .CK (n_121_66), .D (sps__n71));
DFF_X1 \values_reg[53][2]  (.Q (\values[53] [2] ), .CK (n_121_66), .D (spc__n157));
DFF_X1 \values_reg[53][3]  (.Q (\values[53] [3] ), .CK (n_121_66), .D (sps__n78));
DFF_X1 \values_reg[53][4]  (.Q (\values[53] [4] ), .CK (n_121_66), .D (sps__n89));
DFF_X1 \values_reg[53][5]  (.Q (\values[53] [5] ), .CK (n_121_66), .D (spc__n132));
DFF_X1 \values_reg[53][6]  (.Q (\values[53] [6] ), .CK (n_121_66), .D (sps__n118));
DFF_X1 \values_reg[53][7]  (.Q (\values[53] [7] ), .CK (n_121_66), .D (spc__n126));
DFF_X1 \values_reg[53][8]  (.Q (\values[53] [8] ), .CK (n_121_66), .D (sps__n97));
DFF_X1 \values_reg[53][9]  (.Q (\values[53] [9] ), .CK (n_121_66), .D (sps__n109));
DFF_X1 \values_reg[53][10]  (.Q (\values[53] [10] ), .CK (n_121_66), .D (sps__n1));
DFF_X1 \values_reg[53][11]  (.Q (\values[53] [11] ), .CK (n_121_66), .D (sps__n12));
DFF_X1 \values_reg[53][12]  (.Q (\values[53] [12] ), .CK (n_121_66), .D (sps__n55));
DFF_X1 \values_reg[53][13]  (.Q (\values[53] [13] ), .CK (n_121_66), .D (sps__n40));
DFF_X1 \values_reg[53][14]  (.Q (\values[53] [14] ), .CK (n_121_66), .D (sps__n28));
DFF_X1 \values_reg[53][15]  (.Q (\values[53] [15] ), .CK (n_121_66), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[53]_reg  (.GCK (n_121_66), .CK (clk), .E (n_53), .SE (1'b0 ));
DFF_X1 \values_reg[54][0]  (.Q (\values[54] [0] ), .CK (n_121_65), .D (sps__n5));
DFF_X1 \values_reg[54][1]  (.Q (\values[54] [1] ), .CK (n_121_65), .D (sps__n71));
DFF_X1 \values_reg[54][2]  (.Q (\values[54] [2] ), .CK (n_121_65), .D (spc__n158));
DFF_X1 \values_reg[54][3]  (.Q (\values[54] [3] ), .CK (n_121_65), .D (sps__n79));
DFF_X1 \values_reg[54][4]  (.Q (\values[54] [4] ), .CK (n_121_65), .D (sps__n89));
DFF_X1 \values_reg[54][5]  (.Q (\values[54] [5] ), .CK (n_121_65), .D (spc__n132));
DFF_X1 \values_reg[54][6]  (.Q (\values[54] [6] ), .CK (n_121_65), .D (sps__n119));
DFF_X1 \values_reg[54][7]  (.Q (\values[54] [7] ), .CK (n_121_65), .D (spc__n126));
DFF_X1 \values_reg[54][8]  (.Q (\values[54] [8] ), .CK (n_121_65), .D (sps__n97));
DFF_X1 \values_reg[54][9]  (.Q (\values[54] [9] ), .CK (n_121_65), .D (sps__n110));
DFF_X1 \values_reg[54][10]  (.Q (\values[54] [10] ), .CK (n_121_65), .D (sps__n1));
DFF_X1 \values_reg[54][11]  (.Q (\values[54] [11] ), .CK (n_121_65), .D (sps__n14));
DFF_X1 \values_reg[54][12]  (.Q (\values[54] [12] ), .CK (n_121_65), .D (sps__n55));
DFF_X1 \values_reg[54][13]  (.Q (\values[54] [13] ), .CK (n_121_65), .D (sps__n38));
DFF_X1 \values_reg[54][14]  (.Q (\values[54] [14] ), .CK (n_121_65), .D (sps__n28));
DFF_X1 \values_reg[54][15]  (.Q (\values[54] [15] ), .CK (n_121_65), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[54]_reg  (.GCK (n_121_65), .CK (clk), .E (n_54), .SE (1'b0 ));
DFF_X1 \values_reg[55][0]  (.Q (\values[55] [0] ), .CK (n_121_64), .D (sps__n5));
DFF_X1 \values_reg[55][1]  (.Q (\values[55] [1] ), .CK (n_121_64), .D (sps__n71));
DFF_X1 \values_reg[55][2]  (.Q (\values[55] [2] ), .CK (n_121_64), .D (spc__n157));
DFF_X1 \values_reg[55][3]  (.Q (\values[55] [3] ), .CK (n_121_64), .D (sps__n78));
DFF_X1 \values_reg[55][4]  (.Q (\values[55] [4] ), .CK (n_121_64), .D (sps__n89));
DFF_X1 \values_reg[55][5]  (.Q (\values[55] [5] ), .CK (n_121_64), .D (spc__n132));
DFF_X1 \values_reg[55][6]  (.Q (\values[55] [6] ), .CK (n_121_64), .D (sps__n118));
DFF_X1 \values_reg[55][7]  (.Q (\values[55] [7] ), .CK (n_121_64), .D (spc__n126));
DFF_X1 \values_reg[55][8]  (.Q (\values[55] [8] ), .CK (n_121_64), .D (sps__n97));
DFF_X1 \values_reg[55][9]  (.Q (\values[55] [9] ), .CK (n_121_64), .D (sps__n109));
DFF_X1 \values_reg[55][10]  (.Q (\values[55] [10] ), .CK (n_121_64), .D (sps__n1));
DFF_X1 \values_reg[55][11]  (.Q (\values[55] [11] ), .CK (n_121_64), .D (sps__n12));
DFF_X1 \values_reg[55][12]  (.Q (\values[55] [12] ), .CK (n_121_64), .D (sps__n52));
DFF_X1 \values_reg[55][13]  (.Q (\values[55] [13] ), .CK (n_121_64), .D (sps__n40));
DFF_X1 \values_reg[55][14]  (.Q (\values[55] [14] ), .CK (n_121_64), .D (sps__n28));
DFF_X1 \values_reg[55][15]  (.Q (\values[55] [15] ), .CK (n_121_64), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[55]_reg  (.GCK (n_121_64), .CK (clk), .E (n_55), .SE (1'b0 ));
DFF_X1 \values_reg[56][0]  (.Q (\values[56] [0] ), .CK (n_121_63), .D (sps__n5));
DFF_X1 \values_reg[56][1]  (.Q (\values[56] [1] ), .CK (n_121_63), .D (sps__n71));
DFF_X1 \values_reg[56][2]  (.Q (\values[56] [2] ), .CK (n_121_63), .D (spc__n157));
DFF_X1 \values_reg[56][3]  (.Q (\values[56] [3] ), .CK (n_121_63), .D (sps__n79));
DFF_X1 \values_reg[56][4]  (.Q (\values[56] [4] ), .CK (n_121_63), .D (sps__n89));
DFF_X1 \values_reg[56][5]  (.Q (\values[56] [5] ), .CK (n_121_63), .D (spc__n132));
DFF_X1 \values_reg[56][6]  (.Q (\values[56] [6] ), .CK (n_121_63), .D (sps__n118));
DFF_X1 \values_reg[56][7]  (.Q (\values[56] [7] ), .CK (n_121_63), .D (spc__n126));
DFF_X1 \values_reg[56][8]  (.Q (\values[56] [8] ), .CK (n_121_63), .D (sps__n97));
DFF_X1 \values_reg[56][9]  (.Q (\values[56] [9] ), .CK (n_121_63), .D (sps__n109));
DFF_X1 \values_reg[56][10]  (.Q (\values[56] [10] ), .CK (n_121_63), .D (sps__n1));
DFF_X1 \values_reg[56][11]  (.Q (\values[56] [11] ), .CK (n_121_63), .D (sps__n14));
DFF_X1 \values_reg[56][12]  (.Q (\values[56] [12] ), .CK (n_121_63), .D (sps__n55));
DFF_X1 \values_reg[56][13]  (.Q (\values[56] [13] ), .CK (n_121_63), .D (sps__n40));
DFF_X1 \values_reg[56][14]  (.Q (\values[56] [14] ), .CK (n_121_63), .D (sps__n28));
DFF_X1 \values_reg[56][15]  (.Q (\values[56] [15] ), .CK (n_121_63), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[56]_reg  (.GCK (n_121_63), .CK (clk), .E (n_56), .SE (1'b0 ));
DFF_X1 \values_reg[57][0]  (.Q (\values[57] [0] ), .CK (n_121_62), .D (sps__n5));
DFF_X1 \values_reg[57][1]  (.Q (\values[57] [1] ), .CK (n_121_62), .D (sps__n71));
DFF_X1 \values_reg[57][2]  (.Q (\values[57] [2] ), .CK (n_121_62), .D (spc__n157));
DFF_X1 \values_reg[57][3]  (.Q (\values[57] [3] ), .CK (n_121_62), .D (sps__n79));
DFF_X1 \values_reg[57][4]  (.Q (\values[57] [4] ), .CK (n_121_62), .D (sps__n89));
DFF_X1 \values_reg[57][5]  (.Q (\values[57] [5] ), .CK (n_121_62), .D (spc__n132));
DFF_X1 \values_reg[57][6]  (.Q (\values[57] [6] ), .CK (n_121_62), .D (sps__n118));
DFF_X1 \values_reg[57][7]  (.Q (\values[57] [7] ), .CK (n_121_62), .D (spc__n126));
DFF_X1 \values_reg[57][8]  (.Q (\values[57] [8] ), .CK (n_121_62), .D (sps__n97));
DFF_X1 \values_reg[57][9]  (.Q (\values[57] [9] ), .CK (n_121_62), .D (sps__n109));
DFF_X1 \values_reg[57][10]  (.Q (\values[57] [10] ), .CK (n_121_62), .D (sps__n1));
DFF_X1 \values_reg[57][11]  (.Q (\values[57] [11] ), .CK (n_121_62), .D (sps__n14));
DFF_X1 \values_reg[57][12]  (.Q (\values[57] [12] ), .CK (n_121_62), .D (sps__n55));
DFF_X1 \values_reg[57][13]  (.Q (\values[57] [13] ), .CK (n_121_62), .D (sps__n40));
DFF_X1 \values_reg[57][14]  (.Q (\values[57] [14] ), .CK (n_121_62), .D (sps__n28));
DFF_X1 \values_reg[57][15]  (.Q (\values[57] [15] ), .CK (n_121_62), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[57]_reg  (.GCK (n_121_62), .CK (clk), .E (n_57), .SE (1'b0 ));
DFF_X1 \values_reg[58][0]  (.Q (\values[58] [0] ), .CK (n_121_61), .D (sps__n5));
DFF_X1 \values_reg[58][1]  (.Q (\values[58] [1] ), .CK (n_121_61), .D (sps__n71));
DFF_X1 \values_reg[58][2]  (.Q (\values[58] [2] ), .CK (n_121_61), .D (spc__n157));
DFF_X1 \values_reg[58][3]  (.Q (\values[58] [3] ), .CK (n_121_61), .D (sps__n79));
DFF_X1 \values_reg[58][4]  (.Q (\values[58] [4] ), .CK (n_121_61), .D (sps__n89));
DFF_X1 \values_reg[58][5]  (.Q (\values[58] [5] ), .CK (n_121_61), .D (spc__n132));
DFF_X1 \values_reg[58][6]  (.Q (\values[58] [6] ), .CK (n_121_61), .D (sps__n118));
DFF_X1 \values_reg[58][7]  (.Q (\values[58] [7] ), .CK (n_121_61), .D (spc__n126));
DFF_X1 \values_reg[58][8]  (.Q (\values[58] [8] ), .CK (n_121_61), .D (sps__n97));
DFF_X1 \values_reg[58][9]  (.Q (\values[58] [9] ), .CK (n_121_61), .D (sps__n109));
DFF_X1 \values_reg[58][10]  (.Q (\values[58] [10] ), .CK (n_121_61), .D (sps__n1));
DFF_X1 \values_reg[58][11]  (.Q (\values[58] [11] ), .CK (n_121_61), .D (sps__n14));
DFF_X1 \values_reg[58][12]  (.Q (\values[58] [12] ), .CK (n_121_61), .D (sps__n55));
DFF_X1 \values_reg[58][13]  (.Q (\values[58] [13] ), .CK (n_121_61), .D (sps__n40));
DFF_X1 \values_reg[58][14]  (.Q (\values[58] [14] ), .CK (n_121_61), .D (sps__n28));
DFF_X1 \values_reg[58][15]  (.Q (\values[58] [15] ), .CK (n_121_61), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[58]_reg  (.GCK (n_121_61), .CK (clk), .E (n_58), .SE (1'b0 ));
DFF_X1 \values_reg[59][0]  (.Q (\values[59] [0] ), .CK (n_121_60), .D (sps__n5));
DFF_X1 \values_reg[59][1]  (.Q (\values[59] [1] ), .CK (n_121_60), .D (sps__n71));
DFF_X1 \values_reg[59][2]  (.Q (\values[59] [2] ), .CK (n_121_60), .D (spc__n157));
DFF_X1 \values_reg[59][3]  (.Q (\values[59] [3] ), .CK (n_121_60), .D (sps__n79));
DFF_X1 \values_reg[59][4]  (.Q (\values[59] [4] ), .CK (n_121_60), .D (sps__n89));
DFF_X1 \values_reg[59][5]  (.Q (\values[59] [5] ), .CK (n_121_60), .D (spc__n132));
DFF_X1 \values_reg[59][6]  (.Q (\values[59] [6] ), .CK (n_121_60), .D (sps__n118));
DFF_X1 \values_reg[59][7]  (.Q (\values[59] [7] ), .CK (n_121_60), .D (spc__n126));
DFF_X1 \values_reg[59][8]  (.Q (\values[59] [8] ), .CK (n_121_60), .D (sps__n97));
DFF_X1 \values_reg[59][9]  (.Q (\values[59] [9] ), .CK (n_121_60), .D (sps__n109));
DFF_X1 \values_reg[59][10]  (.Q (\values[59] [10] ), .CK (n_121_60), .D (sps__n1));
DFF_X1 \values_reg[59][11]  (.Q (\values[59] [11] ), .CK (n_121_60), .D (sps__n14));
DFF_X1 \values_reg[59][12]  (.Q (\values[59] [12] ), .CK (n_121_60), .D (sps__n55));
DFF_X1 \values_reg[59][13]  (.Q (\values[59] [13] ), .CK (n_121_60), .D (sps__n40));
DFF_X1 \values_reg[59][14]  (.Q (\values[59] [14] ), .CK (n_121_60), .D (sps__n28));
DFF_X1 \values_reg[59][15]  (.Q (\values[59] [15] ), .CK (n_121_60), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[59]_reg  (.GCK (n_121_60), .CK (clk), .E (n_59), .SE (1'b0 ));
DFF_X1 \values_reg[60][0]  (.Q (\values[60] [0] ), .CK (n_121_59), .D (sps__n5));
DFF_X1 \values_reg[60][1]  (.Q (\values[60] [1] ), .CK (n_121_59), .D (sps__n71));
DFF_X1 \values_reg[60][2]  (.Q (\values[60] [2] ), .CK (n_121_59), .D (spc__n157));
DFF_X1 \values_reg[60][3]  (.Q (\values[60] [3] ), .CK (n_121_59), .D (sps__n79));
DFF_X1 \values_reg[60][4]  (.Q (\values[60] [4] ), .CK (n_121_59), .D (sps__n89));
DFF_X1 \values_reg[60][5]  (.Q (\values[60] [5] ), .CK (n_121_59), .D (spc__n132));
DFF_X1 \values_reg[60][6]  (.Q (\values[60] [6] ), .CK (n_121_59), .D (sps__n118));
DFF_X1 \values_reg[60][7]  (.Q (\values[60] [7] ), .CK (n_121_59), .D (spc__n126));
DFF_X1 \values_reg[60][8]  (.Q (\values[60] [8] ), .CK (n_121_59), .D (sps__n97));
DFF_X1 \values_reg[60][9]  (.Q (\values[60] [9] ), .CK (n_121_59), .D (sps__n109));
DFF_X1 \values_reg[60][10]  (.Q (\values[60] [10] ), .CK (n_121_59), .D (sps__n1));
DFF_X1 \values_reg[60][11]  (.Q (\values[60] [11] ), .CK (n_121_59), .D (sps__n14));
DFF_X1 \values_reg[60][12]  (.Q (\values[60] [12] ), .CK (n_121_59), .D (sps__n55));
DFF_X1 \values_reg[60][13]  (.Q (\values[60] [13] ), .CK (n_121_59), .D (sps__n40));
DFF_X1 \values_reg[60][14]  (.Q (\values[60] [14] ), .CK (n_121_59), .D (sps__n28));
DFF_X1 \values_reg[60][15]  (.Q (\values[60] [15] ), .CK (n_121_59), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[60]_reg  (.GCK (n_121_59), .CK (clk), .E (n_60), .SE (1'b0 ));
DFF_X1 \values_reg[61][0]  (.Q (\values[61] [0] ), .CK (n_121_58), .D (sps__n5));
DFF_X1 \values_reg[61][1]  (.Q (\values[61] [1] ), .CK (n_121_58), .D (sps__n71));
DFF_X1 \values_reg[61][2]  (.Q (\values[61] [2] ), .CK (n_121_58), .D (spc__n157));
DFF_X1 \values_reg[61][3]  (.Q (\values[61] [3] ), .CK (n_121_58), .D (sps__n79));
DFF_X1 \values_reg[61][4]  (.Q (\values[61] [4] ), .CK (n_121_58), .D (sps__n89));
DFF_X1 \values_reg[61][5]  (.Q (\values[61] [5] ), .CK (n_121_58), .D (spc__n132));
DFF_X1 \values_reg[61][6]  (.Q (\values[61] [6] ), .CK (n_121_58), .D (sps__n118));
DFF_X1 \values_reg[61][7]  (.Q (\values[61] [7] ), .CK (n_121_58), .D (spc__n126));
DFF_X1 \values_reg[61][8]  (.Q (\values[61] [8] ), .CK (n_121_58), .D (sps__n97));
DFF_X1 \values_reg[61][9]  (.Q (\values[61] [9] ), .CK (n_121_58), .D (sps__n109));
DFF_X1 \values_reg[61][10]  (.Q (\values[61] [10] ), .CK (n_121_58), .D (sps__n1));
DFF_X1 \values_reg[61][11]  (.Q (\values[61] [11] ), .CK (n_121_58), .D (sps__n12));
DFF_X1 \values_reg[61][12]  (.Q (\values[61] [12] ), .CK (n_121_58), .D (sps__n55));
DFF_X1 \values_reg[61][13]  (.Q (\values[61] [13] ), .CK (n_121_58), .D (sps__n40));
DFF_X1 \values_reg[61][14]  (.Q (\values[61] [14] ), .CK (n_121_58), .D (sps__n28));
DFF_X1 \values_reg[61][15]  (.Q (\values[61] [15] ), .CK (n_121_58), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[61]_reg  (.GCK (n_121_58), .CK (clk), .E (n_61), .SE (1'b0 ));
DFF_X1 \values_reg[62][0]  (.Q (\values[62] [0] ), .CK (n_121_57), .D (sps__n5));
DFF_X1 \values_reg[62][1]  (.Q (\values[62] [1] ), .CK (n_121_57), .D (sps__n71));
DFF_X1 \values_reg[62][2]  (.Q (\values[62] [2] ), .CK (n_121_57), .D (spc__n157));
DFF_X1 \values_reg[62][3]  (.Q (\values[62] [3] ), .CK (n_121_57), .D (sps__n79));
DFF_X1 \values_reg[62][4]  (.Q (\values[62] [4] ), .CK (n_121_57), .D (sps__n89));
DFF_X1 \values_reg[62][5]  (.Q (\values[62] [5] ), .CK (n_121_57), .D (spc__n132));
DFF_X1 \values_reg[62][6]  (.Q (\values[62] [6] ), .CK (n_121_57), .D (sps__n118));
DFF_X1 \values_reg[62][7]  (.Q (\values[62] [7] ), .CK (n_121_57), .D (spc__n126));
DFF_X1 \values_reg[62][8]  (.Q (\values[62] [8] ), .CK (n_121_57), .D (sps__n97));
DFF_X1 \values_reg[62][9]  (.Q (\values[62] [9] ), .CK (n_121_57), .D (sps__n109));
DFF_X1 \values_reg[62][10]  (.Q (\values[62] [10] ), .CK (n_121_57), .D (sps__n1));
DFF_X1 \values_reg[62][11]  (.Q (\values[62] [11] ), .CK (n_121_57), .D (sps__n14));
DFF_X1 \values_reg[62][12]  (.Q (\values[62] [12] ), .CK (n_121_57), .D (sps__n55));
DFF_X1 \values_reg[62][13]  (.Q (\values[62] [13] ), .CK (n_121_57), .D (sps__n40));
DFF_X1 \values_reg[62][14]  (.Q (\values[62] [14] ), .CK (n_121_57), .D (sps__n28));
DFF_X1 \values_reg[62][15]  (.Q (\values[62] [15] ), .CK (n_121_57), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[62]_reg  (.GCK (n_121_57), .CK (clk), .E (n_62), .SE (1'b0 ));
DFF_X1 \values_reg[63][0]  (.Q (\values[63] [0] ), .CK (n_121_56), .D (sps__n5));
DFF_X1 \values_reg[63][1]  (.Q (\values[63] [1] ), .CK (n_121_56), .D (sps__n71));
DFF_X1 \values_reg[63][2]  (.Q (\values[63] [2] ), .CK (n_121_56), .D (spc__n157));
DFF_X1 \values_reg[63][3]  (.Q (\values[63] [3] ), .CK (n_121_56), .D (sps__n79));
DFF_X1 \values_reg[63][4]  (.Q (\values[63] [4] ), .CK (n_121_56), .D (sps__n89));
DFF_X1 \values_reg[63][5]  (.Q (\values[63] [5] ), .CK (n_121_56), .D (spc__n132));
DFF_X1 \values_reg[63][6]  (.Q (\values[63] [6] ), .CK (n_121_56), .D (sps__n118));
DFF_X1 \values_reg[63][7]  (.Q (\values[63] [7] ), .CK (n_121_56), .D (spc__n126));
DFF_X1 \values_reg[63][8]  (.Q (\values[63] [8] ), .CK (n_121_56), .D (sps__n97));
DFF_X1 \values_reg[63][9]  (.Q (\values[63] [9] ), .CK (n_121_56), .D (sps__n109));
DFF_X1 \values_reg[63][10]  (.Q (\values[63] [10] ), .CK (n_121_56), .D (sps__n1));
DFF_X1 \values_reg[63][11]  (.Q (\values[63] [11] ), .CK (n_121_56), .D (sps__n12));
DFF_X1 \values_reg[63][12]  (.Q (\values[63] [12] ), .CK (n_121_56), .D (sps__n55));
DFF_X1 \values_reg[63][13]  (.Q (\values[63] [13] ), .CK (n_121_56), .D (sps__n40));
DFF_X1 \values_reg[63][14]  (.Q (\values[63] [14] ), .CK (n_121_56), .D (sps__n28));
DFF_X1 \values_reg[63][15]  (.Q (\values[63] [15] ), .CK (n_121_56), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[63]_reg  (.GCK (n_121_56), .CK (clk), .E (n_63), .SE (1'b0 ));
DFF_X1 \values_reg[64][0]  (.Q (\values[64] [0] ), .CK (n_121_55), .D (sps__n5));
DFF_X1 \values_reg[64][1]  (.Q (\values[64] [1] ), .CK (n_121_55), .D (sps__n71));
DFF_X1 \values_reg[64][2]  (.Q (\values[64] [2] ), .CK (n_121_55), .D (spc__n157));
DFF_X1 \values_reg[64][3]  (.Q (\values[64] [3] ), .CK (n_121_55), .D (sps__n79));
DFF_X1 \values_reg[64][4]  (.Q (\values[64] [4] ), .CK (n_121_55), .D (sps__n89));
DFF_X1 \values_reg[64][5]  (.Q (\values[64] [5] ), .CK (n_121_55), .D (spc__n132));
DFF_X1 \values_reg[64][6]  (.Q (\values[64] [6] ), .CK (n_121_55), .D (sps__n118));
DFF_X1 \values_reg[64][7]  (.Q (\values[64] [7] ), .CK (n_121_55), .D (spc__n126));
DFF_X1 \values_reg[64][8]  (.Q (\values[64] [8] ), .CK (n_121_55), .D (sps__n97));
DFF_X1 \values_reg[64][9]  (.Q (\values[64] [9] ), .CK (n_121_55), .D (sps__n109));
DFF_X1 \values_reg[64][10]  (.Q (\values[64] [10] ), .CK (n_121_55), .D (sps__n1));
DFF_X1 \values_reg[64][11]  (.Q (\values[64] [11] ), .CK (n_121_55), .D (sps__n12));
DFF_X1 \values_reg[64][12]  (.Q (\values[64] [12] ), .CK (n_121_55), .D (sps__n55));
DFF_X1 \values_reg[64][13]  (.Q (\values[64] [13] ), .CK (n_121_55), .D (sps__n40));
DFF_X1 \values_reg[64][14]  (.Q (\values[64] [14] ), .CK (n_121_55), .D (sps__n28));
DFF_X1 \values_reg[64][15]  (.Q (\values[64] [15] ), .CK (n_121_55), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[64]_reg  (.GCK (n_121_55), .CK (clk), .E (n_64), .SE (1'b0 ));
DFF_X1 \values_reg[65][0]  (.Q (\values[65] [0] ), .CK (n_121_54), .D (sps__n5));
DFF_X1 \values_reg[65][1]  (.Q (\values[65] [1] ), .CK (n_121_54), .D (sps__n71));
DFF_X1 \values_reg[65][2]  (.Q (\values[65] [2] ), .CK (n_121_54), .D (spc__n157));
DFF_X1 \values_reg[65][3]  (.Q (\values[65] [3] ), .CK (n_121_54), .D (sps__n79));
DFF_X1 \values_reg[65][4]  (.Q (\values[65] [4] ), .CK (n_121_54), .D (sps__n89));
DFF_X1 \values_reg[65][5]  (.Q (\values[65] [5] ), .CK (n_121_54), .D (spc__n132));
DFF_X1 \values_reg[65][6]  (.Q (\values[65] [6] ), .CK (n_121_54), .D (sps__n118));
DFF_X1 \values_reg[65][7]  (.Q (\values[65] [7] ), .CK (n_121_54), .D (spc__n126));
DFF_X1 \values_reg[65][8]  (.Q (\values[65] [8] ), .CK (n_121_54), .D (sps__n97));
DFF_X1 \values_reg[65][9]  (.Q (\values[65] [9] ), .CK (n_121_54), .D (sps__n109));
DFF_X1 \values_reg[65][10]  (.Q (\values[65] [10] ), .CK (n_121_54), .D (sps__n1));
DFF_X1 \values_reg[65][11]  (.Q (\values[65] [11] ), .CK (n_121_54), .D (sps__n12));
DFF_X1 \values_reg[65][12]  (.Q (\values[65] [12] ), .CK (n_121_54), .D (sps__n55));
DFF_X1 \values_reg[65][13]  (.Q (\values[65] [13] ), .CK (n_121_54), .D (sps__n40));
DFF_X1 \values_reg[65][14]  (.Q (\values[65] [14] ), .CK (n_121_54), .D (sps__n28));
DFF_X1 \values_reg[65][15]  (.Q (\values[65] [15] ), .CK (n_121_54), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[65]_reg  (.GCK (n_121_54), .CK (clk), .E (n_65), .SE (1'b0 ));
DFF_X1 \values_reg[66][0]  (.Q (\values[66] [0] ), .CK (n_121_53), .D (sps__n5));
DFF_X1 \values_reg[66][1]  (.Q (\values[66] [1] ), .CK (n_121_53), .D (sps__n71));
DFF_X1 \values_reg[66][2]  (.Q (\values[66] [2] ), .CK (n_121_53), .D (spc__n159));
DFF_X1 \values_reg[66][3]  (.Q (\values[66] [3] ), .CK (n_121_53), .D (sps__n77));
DFF_X1 \values_reg[66][4]  (.Q (\values[66] [4] ), .CK (n_121_53), .D (sps__n89));
DFF_X1 \values_reg[66][5]  (.Q (\values[66] [5] ), .CK (n_121_53), .D (spc__n132));
DFF_X1 \values_reg[66][6]  (.Q (\values[66] [6] ), .CK (n_121_53), .D (sps__n118));
DFF_X1 \values_reg[66][7]  (.Q (\values[66] [7] ), .CK (n_121_53), .D (spc__n127));
DFF_X1 \values_reg[66][8]  (.Q (\values[66] [8] ), .CK (n_121_53), .D (sps__n97));
DFF_X1 \values_reg[66][9]  (.Q (\values[66] [9] ), .CK (n_121_53), .D (sps__n109));
DFF_X1 \values_reg[66][10]  (.Q (\values[66] [10] ), .CK (n_121_53), .D (sps__n1));
DFF_X1 \values_reg[66][11]  (.Q (\values[66] [11] ), .CK (n_121_53), .D (sps__n12));
DFF_X1 \values_reg[66][12]  (.Q (\values[66] [12] ), .CK (n_121_53), .D (sps__n54));
DFF_X1 \values_reg[66][13]  (.Q (\values[66] [13] ), .CK (n_121_53), .D (sps__n39));
DFF_X1 \values_reg[66][14]  (.Q (\values[66] [14] ), .CK (n_121_53), .D (sps__n27));
DFF_X1 \values_reg[66][15]  (.Q (\values[66] [15] ), .CK (n_121_53), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[66]_reg  (.GCK (n_121_53), .CK (clk), .E (n_66), .SE (1'b0 ));
DFF_X1 \values_reg[67][0]  (.Q (\values[67] [0] ), .CK (n_121_52), .D (sps__n5));
DFF_X1 \values_reg[67][1]  (.Q (\values[67] [1] ), .CK (n_121_52), .D (sps__n71));
DFF_X1 \values_reg[67][2]  (.Q (\values[67] [2] ), .CK (n_121_52), .D (spc__n159));
DFF_X1 \values_reg[67][3]  (.Q (\values[67] [3] ), .CK (n_121_52), .D (sps__n77));
DFF_X1 \values_reg[67][4]  (.Q (\values[67] [4] ), .CK (n_121_52), .D (sps__n89));
DFF_X1 \values_reg[67][5]  (.Q (\values[67] [5] ), .CK (n_121_52), .D (spc__n132));
DFF_X1 \values_reg[67][6]  (.Q (\values[67] [6] ), .CK (n_121_52), .D (sps__n118));
DFF_X1 \values_reg[67][7]  (.Q (\values[67] [7] ), .CK (n_121_52), .D (spc__n127));
DFF_X1 \values_reg[67][8]  (.Q (\values[67] [8] ), .CK (n_121_52), .D (sps__n97));
DFF_X1 \values_reg[67][9]  (.Q (\values[67] [9] ), .CK (n_121_52), .D (sps__n109));
DFF_X1 \values_reg[67][10]  (.Q (\values[67] [10] ), .CK (n_121_52), .D (sps__n1));
DFF_X1 \values_reg[67][11]  (.Q (\values[67] [11] ), .CK (n_121_52), .D (sps__n12));
DFF_X1 \values_reg[67][12]  (.Q (\values[67] [12] ), .CK (n_121_52), .D (sps__n54));
DFF_X1 \values_reg[67][13]  (.Q (\values[67] [13] ), .CK (n_121_52), .D (sps__n40));
DFF_X1 \values_reg[67][14]  (.Q (\values[67] [14] ), .CK (n_121_52), .D (sps__n28));
DFF_X1 \values_reg[67][15]  (.Q (\values[67] [15] ), .CK (n_121_52), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[67]_reg  (.GCK (n_121_52), .CK (clk), .E (n_67), .SE (1'b0 ));
DFF_X1 \values_reg[68][0]  (.Q (\values[68] [0] ), .CK (n_121_51), .D (sps__n5));
DFF_X1 \values_reg[68][1]  (.Q (\values[68] [1] ), .CK (n_121_51), .D (sps__n71));
DFF_X1 \values_reg[68][2]  (.Q (\values[68] [2] ), .CK (n_121_51), .D (spc__n157));
DFF_X1 \values_reg[68][3]  (.Q (\values[68] [3] ), .CK (n_121_51), .D (sps__n79));
DFF_X1 \values_reg[68][4]  (.Q (\values[68] [4] ), .CK (n_121_51), .D (sps__n89));
DFF_X1 \values_reg[68][5]  (.Q (\values[68] [5] ), .CK (n_121_51), .D (spc__n132));
DFF_X1 \values_reg[68][6]  (.Q (\values[68] [6] ), .CK (n_121_51), .D (sps__n118));
DFF_X1 \values_reg[68][7]  (.Q (\values[68] [7] ), .CK (n_121_51), .D (spc__n126));
DFF_X1 \values_reg[68][8]  (.Q (\values[68] [8] ), .CK (n_121_51), .D (sps__n97));
DFF_X1 \values_reg[68][9]  (.Q (\values[68] [9] ), .CK (n_121_51), .D (sps__n110));
DFF_X1 \values_reg[68][10]  (.Q (\values[68] [10] ), .CK (n_121_51), .D (sps__n1));
DFF_X1 \values_reg[68][11]  (.Q (\values[68] [11] ), .CK (n_121_51), .D (sps__n12));
DFF_X1 \values_reg[68][12]  (.Q (\values[68] [12] ), .CK (n_121_51), .D (sps__n55));
DFF_X1 \values_reg[68][13]  (.Q (\values[68] [13] ), .CK (n_121_51), .D (sps__n40));
DFF_X1 \values_reg[68][14]  (.Q (\values[68] [14] ), .CK (n_121_51), .D (sps__n28));
DFF_X1 \values_reg[68][15]  (.Q (\values[68] [15] ), .CK (n_121_51), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[68]_reg  (.GCK (n_121_51), .CK (clk), .E (n_68), .SE (1'b0 ));
DFF_X1 \values_reg[69][0]  (.Q (\values[69] [0] ), .CK (n_121_50), .D (sps__n5));
DFF_X1 \values_reg[69][1]  (.Q (\values[69] [1] ), .CK (n_121_50), .D (sps__n71));
DFF_X1 \values_reg[69][2]  (.Q (\values[69] [2] ), .CK (n_121_50), .D (spc__n157));
DFF_X1 \values_reg[69][3]  (.Q (\values[69] [3] ), .CK (n_121_50), .D (sps__n79));
DFF_X1 \values_reg[69][4]  (.Q (\values[69] [4] ), .CK (n_121_50), .D (sps__n89));
DFF_X1 \values_reg[69][5]  (.Q (\values[69] [5] ), .CK (n_121_50), .D (spc__n132));
DFF_X1 \values_reg[69][6]  (.Q (\values[69] [6] ), .CK (n_121_50), .D (sps__n118));
DFF_X1 \values_reg[69][7]  (.Q (\values[69] [7] ), .CK (n_121_50), .D (spc__n126));
DFF_X1 \values_reg[69][8]  (.Q (\values[69] [8] ), .CK (n_121_50), .D (sps__n97));
DFF_X1 \values_reg[69][9]  (.Q (\values[69] [9] ), .CK (n_121_50), .D (sps__n109));
DFF_X1 \values_reg[69][10]  (.Q (\values[69] [10] ), .CK (n_121_50), .D (sps__n1));
DFF_X1 \values_reg[69][11]  (.Q (\values[69] [11] ), .CK (n_121_50), .D (sps__n12));
DFF_X1 \values_reg[69][12]  (.Q (\values[69] [12] ), .CK (n_121_50), .D (sps__n55));
DFF_X1 \values_reg[69][13]  (.Q (\values[69] [13] ), .CK (n_121_50), .D (sps__n40));
DFF_X1 \values_reg[69][14]  (.Q (\values[69] [14] ), .CK (n_121_50), .D (sps__n28));
DFF_X1 \values_reg[69][15]  (.Q (\values[69] [15] ), .CK (n_121_50), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[69]_reg  (.GCK (n_121_50), .CK (clk), .E (n_69), .SE (1'b0 ));
DFF_X1 \values_reg[70][0]  (.Q (\values[70] [0] ), .CK (n_121_49), .D (sps__n5));
DFF_X1 \values_reg[70][1]  (.Q (\values[70] [1] ), .CK (n_121_49), .D (sps__n71));
DFF_X1 \values_reg[70][2]  (.Q (\values[70] [2] ), .CK (n_121_49), .D (spc__n159));
DFF_X1 \values_reg[70][3]  (.Q (\values[70] [3] ), .CK (n_121_49), .D (sps__n77));
DFF_X1 \values_reg[70][4]  (.Q (\values[70] [4] ), .CK (n_121_49), .D (sps__n89));
DFF_X1 \values_reg[70][5]  (.Q (\values[70] [5] ), .CK (n_121_49), .D (spc__n132));
DFF_X1 \values_reg[70][6]  (.Q (\values[70] [6] ), .CK (n_121_49), .D (sps__n118));
DFF_X1 \values_reg[70][7]  (.Q (\values[70] [7] ), .CK (n_121_49), .D (spc__n127));
DFF_X1 \values_reg[70][8]  (.Q (\values[70] [8] ), .CK (n_121_49), .D (sps__n97));
DFF_X1 \values_reg[70][9]  (.Q (\values[70] [9] ), .CK (n_121_49), .D (sps__n109));
DFF_X1 \values_reg[70][10]  (.Q (\values[70] [10] ), .CK (n_121_49), .D (sps__n1));
DFF_X1 \values_reg[70][11]  (.Q (\values[70] [11] ), .CK (n_121_49), .D (sps__n12));
DFF_X1 \values_reg[70][12]  (.Q (\values[70] [12] ), .CK (n_121_49), .D (sps__n54));
DFF_X1 \values_reg[70][13]  (.Q (\values[70] [13] ), .CK (n_121_49), .D (sps__n40));
DFF_X1 \values_reg[70][14]  (.Q (\values[70] [14] ), .CK (n_121_49), .D (sps__n28));
DFF_X1 \values_reg[70][15]  (.Q (\values[70] [15] ), .CK (n_121_49), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[70]_reg  (.GCK (n_121_49), .CK (clk), .E (n_70), .SE (1'b0 ));
DFF_X1 \values_reg[71][0]  (.Q (\values[71] [0] ), .CK (n_121_48), .D (sps__n5));
DFF_X1 \values_reg[71][1]  (.Q (\values[71] [1] ), .CK (n_121_48), .D (sps__n71));
DFF_X1 \values_reg[71][2]  (.Q (\values[71] [2] ), .CK (n_121_48), .D (spc__n159));
DFF_X1 \values_reg[71][3]  (.Q (\values[71] [3] ), .CK (n_121_48), .D (sps__n77));
DFF_X1 \values_reg[71][4]  (.Q (\values[71] [4] ), .CK (n_121_48), .D (sps__n89));
DFF_X1 \values_reg[71][5]  (.Q (\values[71] [5] ), .CK (n_121_48), .D (spc__n132));
DFF_X1 \values_reg[71][6]  (.Q (\values[71] [6] ), .CK (n_121_48), .D (sps__n118));
DFF_X1 \values_reg[71][7]  (.Q (\values[71] [7] ), .CK (n_121_48), .D (spc__n127));
DFF_X1 \values_reg[71][8]  (.Q (\values[71] [8] ), .CK (n_121_48), .D (sps__n97));
DFF_X1 \values_reg[71][9]  (.Q (\values[71] [9] ), .CK (n_121_48), .D (sps__n109));
DFF_X1 \values_reg[71][10]  (.Q (\values[71] [10] ), .CK (n_121_48), .D (sps__n1));
DFF_X1 \values_reg[71][11]  (.Q (\values[71] [11] ), .CK (n_121_48), .D (sps__n12));
DFF_X1 \values_reg[71][12]  (.Q (\values[71] [12] ), .CK (n_121_48), .D (sps__n54));
DFF_X1 \values_reg[71][13]  (.Q (\values[71] [13] ), .CK (n_121_48), .D (sps__n40));
DFF_X1 \values_reg[71][14]  (.Q (\values[71] [14] ), .CK (n_121_48), .D (sps__n28));
DFF_X1 \values_reg[71][15]  (.Q (\values[71] [15] ), .CK (n_121_48), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[71]_reg  (.GCK (n_121_48), .CK (clk), .E (n_71), .SE (1'b0 ));
DFF_X1 \values_reg[72][0]  (.Q (\values[72] [0] ), .CK (n_121_47), .D (sps__n5));
DFF_X1 \values_reg[72][1]  (.Q (\values[72] [1] ), .CK (n_121_47), .D (sps__n71));
DFF_X1 \values_reg[72][2]  (.Q (\values[72] [2] ), .CK (n_121_47), .D (spc__n159));
DFF_X1 \values_reg[72][3]  (.Q (\values[72] [3] ), .CK (n_121_47), .D (sps__n77));
DFF_X1 \values_reg[72][4]  (.Q (\values[72] [4] ), .CK (n_121_47), .D (sps__n89));
DFF_X1 \values_reg[72][5]  (.Q (\values[72] [5] ), .CK (n_121_47), .D (spc__n132));
DFF_X1 \values_reg[72][6]  (.Q (\values[72] [6] ), .CK (n_121_47), .D (sps__n117));
DFF_X1 \values_reg[72][7]  (.Q (\values[72] [7] ), .CK (n_121_47), .D (spc__n127));
DFF_X1 \values_reg[72][8]  (.Q (\values[72] [8] ), .CK (n_121_47), .D (sps__n97));
DFF_X1 \values_reg[72][9]  (.Q (\values[72] [9] ), .CK (n_121_47), .D (sps__n109));
DFF_X1 \values_reg[72][10]  (.Q (\values[72] [10] ), .CK (n_121_47), .D (sps__n1));
DFF_X1 \values_reg[72][11]  (.Q (\values[72] [11] ), .CK (n_121_47), .D (sps__n12));
DFF_X1 \values_reg[72][12]  (.Q (\values[72] [12] ), .CK (n_121_47), .D (sps__n54));
DFF_X1 \values_reg[72][13]  (.Q (\values[72] [13] ), .CK (n_121_47), .D (sps__n40));
DFF_X1 \values_reg[72][14]  (.Q (\values[72] [14] ), .CK (n_121_47), .D (sps__n25));
DFF_X1 \values_reg[72][15]  (.Q (\values[72] [15] ), .CK (n_121_47), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[72]_reg  (.GCK (n_121_47), .CK (clk), .E (n_72), .SE (1'b0 ));
DFF_X1 \values_reg[73][0]  (.Q (\values[73] [0] ), .CK (n_121_46), .D (sps__n5));
DFF_X1 \values_reg[73][1]  (.Q (\values[73] [1] ), .CK (n_121_46), .D (sps__n71));
DFF_X1 \values_reg[73][2]  (.Q (\values[73] [2] ), .CK (n_121_46), .D (spc__n159));
DFF_X1 \values_reg[73][3]  (.Q (\values[73] [3] ), .CK (n_121_46), .D (sps__n77));
DFF_X1 \values_reg[73][4]  (.Q (\values[73] [4] ), .CK (n_121_46), .D (sps__n89));
DFF_X1 \values_reg[73][5]  (.Q (\values[73] [5] ), .CK (n_121_46), .D (spc__n132));
DFF_X1 \values_reg[73][6]  (.Q (\values[73] [6] ), .CK (n_121_46), .D (sps__n117));
DFF_X1 \values_reg[73][7]  (.Q (\values[73] [7] ), .CK (n_121_46), .D (spc__n127));
DFF_X1 \values_reg[73][8]  (.Q (\values[73] [8] ), .CK (n_121_46), .D (sps__n97));
DFF_X1 \values_reg[73][9]  (.Q (\values[73] [9] ), .CK (n_121_46), .D (sps__n109));
DFF_X1 \values_reg[73][10]  (.Q (\values[73] [10] ), .CK (n_121_46), .D (sps__n1));
DFF_X1 \values_reg[73][11]  (.Q (\values[73] [11] ), .CK (n_121_46), .D (sps__n12));
DFF_X1 \values_reg[73][12]  (.Q (\values[73] [12] ), .CK (n_121_46), .D (sps__n54));
DFF_X1 \values_reg[73][13]  (.Q (\values[73] [13] ), .CK (n_121_46), .D (sps__n40));
DFF_X1 \values_reg[73][14]  (.Q (\values[73] [14] ), .CK (n_121_46), .D (sps__n25));
DFF_X1 \values_reg[73][15]  (.Q (\values[73] [15] ), .CK (n_121_46), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[73]_reg  (.GCK (n_121_46), .CK (clk), .E (n_73), .SE (1'b0 ));
DFF_X1 \values_reg[74][0]  (.Q (\values[74] [0] ), .CK (n_121_45), .D (sps__n5));
DFF_X1 \values_reg[74][1]  (.Q (\values[74] [1] ), .CK (n_121_45), .D (sps__n71));
DFF_X1 \values_reg[74][2]  (.Q (\values[74] [2] ), .CK (n_121_45), .D (spc__n157));
DFF_X1 \values_reg[74][3]  (.Q (\values[74] [3] ), .CK (n_121_45), .D (sps__n79));
DFF_X1 \values_reg[74][4]  (.Q (\values[74] [4] ), .CK (n_121_45), .D (sps__n89));
DFF_X1 \values_reg[74][5]  (.Q (\values[74] [5] ), .CK (n_121_45), .D (spc__n132));
DFF_X1 \values_reg[74][6]  (.Q (\values[74] [6] ), .CK (n_121_45), .D (sps__n118));
DFF_X1 \values_reg[74][7]  (.Q (\values[74] [7] ), .CK (n_121_45), .D (spc__n126));
DFF_X1 \values_reg[74][8]  (.Q (\values[74] [8] ), .CK (n_121_45), .D (sps__n97));
DFF_X1 \values_reg[74][9]  (.Q (\values[74] [9] ), .CK (n_121_45), .D (sps__n109));
DFF_X1 \values_reg[74][10]  (.Q (\values[74] [10] ), .CK (n_121_45), .D (sps__n1));
DFF_X1 \values_reg[74][11]  (.Q (\values[74] [11] ), .CK (n_121_45), .D (sps__n12));
DFF_X1 \values_reg[74][12]  (.Q (\values[74] [12] ), .CK (n_121_45), .D (sps__n55));
DFF_X1 \values_reg[74][13]  (.Q (\values[74] [13] ), .CK (n_121_45), .D (sps__n40));
DFF_X1 \values_reg[74][14]  (.Q (\values[74] [14] ), .CK (n_121_45), .D (sps__n28));
DFF_X1 \values_reg[74][15]  (.Q (\values[74] [15] ), .CK (n_121_45), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[74]_reg  (.GCK (n_121_45), .CK (clk), .E (n_74), .SE (1'b0 ));
DFF_X1 \values_reg[75][0]  (.Q (\values[75] [0] ), .CK (n_121_44), .D (sps__n5));
DFF_X1 \values_reg[75][1]  (.Q (\values[75] [1] ), .CK (n_121_44), .D (sps__n71));
DFF_X1 \values_reg[75][2]  (.Q (\values[75] [2] ), .CK (n_121_44), .D (spc__n157));
DFF_X1 \values_reg[75][3]  (.Q (\values[75] [3] ), .CK (n_121_44), .D (sps__n79));
DFF_X1 \values_reg[75][4]  (.Q (\values[75] [4] ), .CK (n_121_44), .D (sps__n89));
DFF_X1 \values_reg[75][5]  (.Q (\values[75] [5] ), .CK (n_121_44), .D (spc__n132));
DFF_X1 \values_reg[75][6]  (.Q (\values[75] [6] ), .CK (n_121_44), .D (sps__n118));
DFF_X1 \values_reg[75][7]  (.Q (\values[75] [7] ), .CK (n_121_44), .D (spc__n126));
DFF_X1 \values_reg[75][8]  (.Q (\values[75] [8] ), .CK (n_121_44), .D (sps__n97));
DFF_X1 \values_reg[75][9]  (.Q (\values[75] [9] ), .CK (n_121_44), .D (sps__n109));
DFF_X1 \values_reg[75][10]  (.Q (\values[75] [10] ), .CK (n_121_44), .D (sps__n1));
DFF_X1 \values_reg[75][11]  (.Q (\values[75] [11] ), .CK (n_121_44), .D (sps__n12));
DFF_X1 \values_reg[75][12]  (.Q (\values[75] [12] ), .CK (n_121_44), .D (sps__n55));
DFF_X1 \values_reg[75][13]  (.Q (\values[75] [13] ), .CK (n_121_44), .D (sps__n40));
DFF_X1 \values_reg[75][14]  (.Q (\values[75] [14] ), .CK (n_121_44), .D (sps__n28));
DFF_X1 \values_reg[75][15]  (.Q (\values[75] [15] ), .CK (n_121_44), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[75]_reg  (.GCK (n_121_44), .CK (clk), .E (n_75), .SE (1'b0 ));
DFF_X1 \values_reg[76][0]  (.Q (\values[76] [0] ), .CK (n_121_43), .D (sps__n5));
DFF_X1 \values_reg[76][1]  (.Q (\values[76] [1] ), .CK (n_121_43), .D (sps__n71));
DFF_X1 \values_reg[76][2]  (.Q (\values[76] [2] ), .CK (n_121_43), .D (spc__n159));
DFF_X1 \values_reg[76][3]  (.Q (\values[76] [3] ), .CK (n_121_43), .D (sps__n77));
DFF_X1 \values_reg[76][4]  (.Q (\values[76] [4] ), .CK (n_121_43), .D (sps__n89));
DFF_X1 \values_reg[76][5]  (.Q (\values[76] [5] ), .CK (n_121_43), .D (spc__n132));
DFF_X1 \values_reg[76][6]  (.Q (\values[76] [6] ), .CK (n_121_43), .D (sps__n117));
DFF_X1 \values_reg[76][7]  (.Q (\values[76] [7] ), .CK (n_121_43), .D (spc__n127));
DFF_X1 \values_reg[76][8]  (.Q (\values[76] [8] ), .CK (n_121_43), .D (sps__n97));
DFF_X1 \values_reg[76][9]  (.Q (\values[76] [9] ), .CK (n_121_43), .D (sps__n109));
DFF_X1 \values_reg[76][10]  (.Q (\values[76] [10] ), .CK (n_121_43), .D (sps__n1));
DFF_X1 \values_reg[76][11]  (.Q (\values[76] [11] ), .CK (n_121_43), .D (sps__n12));
DFF_X1 \values_reg[76][12]  (.Q (\values[76] [12] ), .CK (n_121_43), .D (sps__n54));
DFF_X1 \values_reg[76][13]  (.Q (\values[76] [13] ), .CK (n_121_43), .D (sps__n40));
DFF_X1 \values_reg[76][14]  (.Q (\values[76] [14] ), .CK (n_121_43), .D (sps__n25));
DFF_X1 \values_reg[76][15]  (.Q (\values[76] [15] ), .CK (n_121_43), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[76]_reg  (.GCK (n_121_43), .CK (clk), .E (n_76), .SE (1'b0 ));
DFF_X1 \values_reg[77][0]  (.Q (\values[77] [0] ), .CK (n_121_42), .D (sps__n5));
DFF_X1 \values_reg[77][1]  (.Q (\values[77] [1] ), .CK (n_121_42), .D (sps__n71));
DFF_X1 \values_reg[77][2]  (.Q (\values[77] [2] ), .CK (n_121_42), .D (spc__n159));
DFF_X1 \values_reg[77][3]  (.Q (\values[77] [3] ), .CK (n_121_42), .D (sps__n77));
DFF_X1 \values_reg[77][4]  (.Q (\values[77] [4] ), .CK (n_121_42), .D (sps__n89));
DFF_X1 \values_reg[77][5]  (.Q (\values[77] [5] ), .CK (n_121_42), .D (spc__n132));
DFF_X1 \values_reg[77][6]  (.Q (\values[77] [6] ), .CK (n_121_42), .D (sps__n117));
DFF_X1 \values_reg[77][7]  (.Q (\values[77] [7] ), .CK (n_121_42), .D (spc__n127));
DFF_X1 \values_reg[77][8]  (.Q (\values[77] [8] ), .CK (n_121_42), .D (sps__n97));
DFF_X1 \values_reg[77][9]  (.Q (\values[77] [9] ), .CK (n_121_42), .D (sps__n109));
DFF_X1 \values_reg[77][10]  (.Q (\values[77] [10] ), .CK (n_121_42), .D (sps__n1));
DFF_X1 \values_reg[77][11]  (.Q (\values[77] [11] ), .CK (n_121_42), .D (sps__n12));
DFF_X1 \values_reg[77][12]  (.Q (\values[77] [12] ), .CK (n_121_42), .D (sps__n54));
DFF_X1 \values_reg[77][13]  (.Q (\values[77] [13] ), .CK (n_121_42), .D (sps__n40));
DFF_X1 \values_reg[77][14]  (.Q (\values[77] [14] ), .CK (n_121_42), .D (sps__n25));
DFF_X1 \values_reg[77][15]  (.Q (\values[77] [15] ), .CK (n_121_42), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[77]_reg  (.GCK (n_121_42), .CK (clk), .E (n_77), .SE (1'b0 ));
DFF_X1 \values_reg[78][0]  (.Q (\values[78] [0] ), .CK (n_121_41), .D (sps__n5));
DFF_X1 \values_reg[78][1]  (.Q (\values[78] [1] ), .CK (n_121_41), .D (sps__n71));
DFF_X1 \values_reg[78][2]  (.Q (\values[78] [2] ), .CK (n_121_41), .D (spc__n157));
DFF_X1 \values_reg[78][3]  (.Q (\values[78] [3] ), .CK (n_121_41), .D (sps__n79));
DFF_X1 \values_reg[78][4]  (.Q (\values[78] [4] ), .CK (n_121_41), .D (sps__n89));
DFF_X1 \values_reg[78][5]  (.Q (\values[78] [5] ), .CK (n_121_41), .D (spc__n132));
DFF_X1 \values_reg[78][6]  (.Q (\values[78] [6] ), .CK (n_121_41), .D (sps__n118));
DFF_X1 \values_reg[78][7]  (.Q (\values[78] [7] ), .CK (n_121_41), .D (spc__n126));
DFF_X1 \values_reg[78][8]  (.Q (\values[78] [8] ), .CK (n_121_41), .D (sps__n97));
DFF_X1 \values_reg[78][9]  (.Q (\values[78] [9] ), .CK (n_121_41), .D (sps__n109));
DFF_X1 \values_reg[78][10]  (.Q (\values[78] [10] ), .CK (n_121_41), .D (sps__n1));
DFF_X1 \values_reg[78][11]  (.Q (\values[78] [11] ), .CK (n_121_41), .D (sps__n12));
DFF_X1 \values_reg[78][12]  (.Q (\values[78] [12] ), .CK (n_121_41), .D (sps__n55));
DFF_X1 \values_reg[78][13]  (.Q (\values[78] [13] ), .CK (n_121_41), .D (sps__n40));
DFF_X1 \values_reg[78][14]  (.Q (\values[78] [14] ), .CK (n_121_41), .D (sps__n28));
DFF_X1 \values_reg[78][15]  (.Q (\values[78] [15] ), .CK (n_121_41), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[78]_reg  (.GCK (n_121_41), .CK (clk), .E (n_78), .SE (1'b0 ));
DFF_X1 \values_reg[79][0]  (.Q (\values[79] [0] ), .CK (n_121_40), .D (sps__n5));
DFF_X1 \values_reg[79][1]  (.Q (\values[79] [1] ), .CK (n_121_40), .D (sps__n71));
DFF_X1 \values_reg[79][2]  (.Q (\values[79] [2] ), .CK (n_121_40), .D (spc__n157));
DFF_X1 \values_reg[79][3]  (.Q (\values[79] [3] ), .CK (n_121_40), .D (sps__n79));
DFF_X1 \values_reg[79][4]  (.Q (\values[79] [4] ), .CK (n_121_40), .D (sps__n89));
DFF_X1 \values_reg[79][5]  (.Q (\values[79] [5] ), .CK (n_121_40), .D (spc__n132));
DFF_X1 \values_reg[79][6]  (.Q (\values[79] [6] ), .CK (n_121_40), .D (sps__n118));
DFF_X1 \values_reg[79][7]  (.Q (\values[79] [7] ), .CK (n_121_40), .D (spc__n126));
DFF_X1 \values_reg[79][8]  (.Q (\values[79] [8] ), .CK (n_121_40), .D (sps__n97));
DFF_X1 \values_reg[79][9]  (.Q (\values[79] [9] ), .CK (n_121_40), .D (sps__n109));
DFF_X1 \values_reg[79][10]  (.Q (\values[79] [10] ), .CK (n_121_40), .D (sps__n1));
DFF_X1 \values_reg[79][11]  (.Q (\values[79] [11] ), .CK (n_121_40), .D (sps__n12));
DFF_X1 \values_reg[79][12]  (.Q (\values[79] [12] ), .CK (n_121_40), .D (sps__n55));
DFF_X1 \values_reg[79][13]  (.Q (\values[79] [13] ), .CK (n_121_40), .D (sps__n40));
DFF_X1 \values_reg[79][14]  (.Q (\values[79] [14] ), .CK (n_121_40), .D (sps__n28));
DFF_X1 \values_reg[79][15]  (.Q (\values[79] [15] ), .CK (n_121_40), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[79]_reg  (.GCK (n_121_40), .CK (clk), .E (n_79), .SE (1'b0 ));
DFF_X1 \values_reg[80][0]  (.Q (\values[80] [0] ), .CK (n_121_39), .D (sps__n5));
DFF_X1 \values_reg[80][1]  (.Q (\values[80] [1] ), .CK (n_121_39), .D (sps__n71));
DFF_X1 \values_reg[80][2]  (.Q (\values[80] [2] ), .CK (n_121_39), .D (spc__n157));
DFF_X1 \values_reg[80][3]  (.Q (\values[80] [3] ), .CK (n_121_39), .D (sps__n79));
DFF_X1 \values_reg[80][4]  (.Q (\values[80] [4] ), .CK (n_121_39), .D (sps__n89));
DFF_X1 \values_reg[80][5]  (.Q (\values[80] [5] ), .CK (n_121_39), .D (spc__n132));
DFF_X1 \values_reg[80][6]  (.Q (\values[80] [6] ), .CK (n_121_39), .D (sps__n118));
DFF_X1 \values_reg[80][7]  (.Q (\values[80] [7] ), .CK (n_121_39), .D (spc__n126));
DFF_X1 \values_reg[80][8]  (.Q (\values[80] [8] ), .CK (n_121_39), .D (sps__n97));
DFF_X1 \values_reg[80][9]  (.Q (\values[80] [9] ), .CK (n_121_39), .D (sps__n109));
DFF_X1 \values_reg[80][10]  (.Q (\values[80] [10] ), .CK (n_121_39), .D (sps__n1));
DFF_X1 \values_reg[80][11]  (.Q (\values[80] [11] ), .CK (n_121_39), .D (sps__n12));
DFF_X1 \values_reg[80][12]  (.Q (\values[80] [12] ), .CK (n_121_39), .D (sps__n55));
DFF_X1 \values_reg[80][13]  (.Q (\values[80] [13] ), .CK (n_121_39), .D (sps__n40));
DFF_X1 \values_reg[80][14]  (.Q (\values[80] [14] ), .CK (n_121_39), .D (sps__n28));
DFF_X1 \values_reg[80][15]  (.Q (\values[80] [15] ), .CK (n_121_39), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[80]_reg  (.GCK (n_121_39), .CK (clk), .E (n_80), .SE (1'b0 ));
DFF_X1 \values_reg[81][0]  (.Q (\values[81] [0] ), .CK (n_121_38), .D (sps__n5));
DFF_X1 \values_reg[81][1]  (.Q (\values[81] [1] ), .CK (n_121_38), .D (sps__n71));
DFF_X1 \values_reg[81][2]  (.Q (\values[81] [2] ), .CK (n_121_38), .D (spc__n157));
DFF_X1 \values_reg[81][3]  (.Q (\values[81] [3] ), .CK (n_121_38), .D (sps__n79));
DFF_X1 \values_reg[81][4]  (.Q (\values[81] [4] ), .CK (n_121_38), .D (sps__n89));
DFF_X1 \values_reg[81][5]  (.Q (\values[81] [5] ), .CK (n_121_38), .D (spc__n132));
DFF_X1 \values_reg[81][6]  (.Q (\values[81] [6] ), .CK (n_121_38), .D (sps__n118));
DFF_X1 \values_reg[81][7]  (.Q (\values[81] [7] ), .CK (n_121_38), .D (spc__n126));
DFF_X1 \values_reg[81][8]  (.Q (\values[81] [8] ), .CK (n_121_38), .D (sps__n97));
DFF_X1 \values_reg[81][9]  (.Q (\values[81] [9] ), .CK (n_121_38), .D (sps__n109));
DFF_X1 \values_reg[81][10]  (.Q (\values[81] [10] ), .CK (n_121_38), .D (sps__n1));
DFF_X1 \values_reg[81][11]  (.Q (\values[81] [11] ), .CK (n_121_38), .D (sps__n12));
DFF_X1 \values_reg[81][12]  (.Q (\values[81] [12] ), .CK (n_121_38), .D (sps__n55));
DFF_X1 \values_reg[81][13]  (.Q (\values[81] [13] ), .CK (n_121_38), .D (sps__n40));
DFF_X1 \values_reg[81][14]  (.Q (\values[81] [14] ), .CK (n_121_38), .D (sps__n28));
DFF_X1 \values_reg[81][15]  (.Q (\values[81] [15] ), .CK (n_121_38), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[81]_reg  (.GCK (n_121_38), .CK (clk), .E (n_81), .SE (1'b0 ));
DFF_X1 \values_reg[82][0]  (.Q (\values[82] [0] ), .CK (n_121_37), .D (sps__n5));
DFF_X1 \values_reg[82][1]  (.Q (\values[82] [1] ), .CK (n_121_37), .D (sps__n71));
DFF_X1 \values_reg[82][2]  (.Q (\values[82] [2] ), .CK (n_121_37), .D (spc__n159));
DFF_X1 \values_reg[82][3]  (.Q (\values[82] [3] ), .CK (n_121_37), .D (sps__n78));
DFF_X1 \values_reg[82][4]  (.Q (\values[82] [4] ), .CK (n_121_37), .D (sps__n89));
DFF_X1 \values_reg[82][5]  (.Q (\values[82] [5] ), .CK (n_121_37), .D (spc__n132));
DFF_X1 \values_reg[82][6]  (.Q (\values[82] [6] ), .CK (n_121_37), .D (sps__n118));
DFF_X1 \values_reg[82][7]  (.Q (\values[82] [7] ), .CK (n_121_37), .D (spc__n127));
DFF_X1 \values_reg[82][8]  (.Q (\values[82] [8] ), .CK (n_121_37), .D (sps__n97));
DFF_X1 \values_reg[82][9]  (.Q (\values[82] [9] ), .CK (n_121_37), .D (sps__n109));
DFF_X1 \values_reg[82][10]  (.Q (\values[82] [10] ), .CK (n_121_37), .D (sps__n1));
DFF_X1 \values_reg[82][11]  (.Q (\values[82] [11] ), .CK (n_121_37), .D (sps__n12));
DFF_X1 \values_reg[82][12]  (.Q (\values[82] [12] ), .CK (n_121_37), .D (sps__n54));
DFF_X1 \values_reg[82][13]  (.Q (\values[82] [13] ), .CK (n_121_37), .D (sps__n40));
DFF_X1 \values_reg[82][14]  (.Q (\values[82] [14] ), .CK (n_121_37), .D (sps__n28));
DFF_X1 \values_reg[82][15]  (.Q (\values[82] [15] ), .CK (n_121_37), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[82]_reg  (.GCK (n_121_37), .CK (clk), .E (n_82), .SE (1'b0 ));
DFF_X1 \values_reg[83][0]  (.Q (\values[83] [0] ), .CK (n_121_36), .D (sps__n5));
DFF_X1 \values_reg[83][1]  (.Q (\values[83] [1] ), .CK (n_121_36), .D (sps__n71));
DFF_X1 \values_reg[83][2]  (.Q (\values[83] [2] ), .CK (n_121_36), .D (spc__n159));
DFF_X1 \values_reg[83][3]  (.Q (\values[83] [3] ), .CK (n_121_36), .D (sps__n78));
DFF_X1 \values_reg[83][4]  (.Q (\values[83] [4] ), .CK (n_121_36), .D (sps__n89));
DFF_X1 \values_reg[83][5]  (.Q (\values[83] [5] ), .CK (n_121_36), .D (spc__n132));
DFF_X1 \values_reg[83][6]  (.Q (\values[83] [6] ), .CK (n_121_36), .D (sps__n118));
DFF_X1 \values_reg[83][7]  (.Q (\values[83] [7] ), .CK (n_121_36), .D (spc__n127));
DFF_X1 \values_reg[83][8]  (.Q (\values[83] [8] ), .CK (n_121_36), .D (sps__n97));
DFF_X1 \values_reg[83][9]  (.Q (\values[83] [9] ), .CK (n_121_36), .D (sps__n109));
DFF_X1 \values_reg[83][10]  (.Q (\values[83] [10] ), .CK (n_121_36), .D (sps__n1));
DFF_X1 \values_reg[83][11]  (.Q (\values[83] [11] ), .CK (n_121_36), .D (sps__n12));
DFF_X1 \values_reg[83][12]  (.Q (\values[83] [12] ), .CK (n_121_36), .D (sps__n54));
DFF_X1 \values_reg[83][13]  (.Q (\values[83] [13] ), .CK (n_121_36), .D (sps__n40));
DFF_X1 \values_reg[83][14]  (.Q (\values[83] [14] ), .CK (n_121_36), .D (sps__n28));
DFF_X1 \values_reg[83][15]  (.Q (\values[83] [15] ), .CK (n_121_36), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[83]_reg  (.GCK (n_121_36), .CK (clk), .E (n_83), .SE (1'b0 ));
DFF_X1 \values_reg[84][0]  (.Q (\values[84] [0] ), .CK (n_121_35), .D (sps__n5));
DFF_X1 \values_reg[84][1]  (.Q (\values[84] [1] ), .CK (n_121_35), .D (sps__n71));
DFF_X1 \values_reg[84][2]  (.Q (\values[84] [2] ), .CK (n_121_35), .D (spc__n157));
DFF_X1 \values_reg[84][3]  (.Q (\values[84] [3] ), .CK (n_121_35), .D (sps__n79));
DFF_X1 \values_reg[84][4]  (.Q (\values[84] [4] ), .CK (n_121_35), .D (sps__n89));
DFF_X1 \values_reg[84][5]  (.Q (\values[84] [5] ), .CK (n_121_35), .D (spc__n132));
DFF_X1 \values_reg[84][6]  (.Q (\values[84] [6] ), .CK (n_121_35), .D (sps__n118));
DFF_X1 \values_reg[84][7]  (.Q (\values[84] [7] ), .CK (n_121_35), .D (spc__n126));
DFF_X1 \values_reg[84][8]  (.Q (\values[84] [8] ), .CK (n_121_35), .D (sps__n97));
DFF_X1 \values_reg[84][9]  (.Q (\values[84] [9] ), .CK (n_121_35), .D (sps__n109));
DFF_X1 \values_reg[84][10]  (.Q (\values[84] [10] ), .CK (n_121_35), .D (sps__n1));
DFF_X1 \values_reg[84][11]  (.Q (\values[84] [11] ), .CK (n_121_35), .D (sps__n12));
DFF_X1 \values_reg[84][12]  (.Q (\values[84] [12] ), .CK (n_121_35), .D (sps__n55));
DFF_X1 \values_reg[84][13]  (.Q (\values[84] [13] ), .CK (n_121_35), .D (sps__n40));
DFF_X1 \values_reg[84][14]  (.Q (\values[84] [14] ), .CK (n_121_35), .D (sps__n28));
DFF_X1 \values_reg[84][15]  (.Q (\values[84] [15] ), .CK (n_121_35), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[84]_reg  (.GCK (n_121_35), .CK (clk), .E (n_84), .SE (1'b0 ));
DFF_X1 \values_reg[85][0]  (.Q (\values[85] [0] ), .CK (n_121_34), .D (sps__n5));
DFF_X1 \values_reg[85][1]  (.Q (\values[85] [1] ), .CK (n_121_34), .D (sps__n71));
DFF_X1 \values_reg[85][2]  (.Q (\values[85] [2] ), .CK (n_121_34), .D (spc__n157));
DFF_X1 \values_reg[85][3]  (.Q (\values[85] [3] ), .CK (n_121_34), .D (sps__n79));
DFF_X1 \values_reg[85][4]  (.Q (\values[85] [4] ), .CK (n_121_34), .D (sps__n89));
DFF_X1 \values_reg[85][5]  (.Q (\values[85] [5] ), .CK (n_121_34), .D (spc__n132));
DFF_X1 \values_reg[85][6]  (.Q (\values[85] [6] ), .CK (n_121_34), .D (sps__n118));
DFF_X1 \values_reg[85][7]  (.Q (\values[85] [7] ), .CK (n_121_34), .D (spc__n126));
DFF_X1 \values_reg[85][8]  (.Q (\values[85] [8] ), .CK (n_121_34), .D (sps__n97));
DFF_X1 \values_reg[85][9]  (.Q (\values[85] [9] ), .CK (n_121_34), .D (sps__n109));
DFF_X1 \values_reg[85][10]  (.Q (\values[85] [10] ), .CK (n_121_34), .D (sps__n1));
DFF_X1 \values_reg[85][11]  (.Q (\values[85] [11] ), .CK (n_121_34), .D (sps__n12));
DFF_X1 \values_reg[85][12]  (.Q (\values[85] [12] ), .CK (n_121_34), .D (sps__n55));
DFF_X1 \values_reg[85][13]  (.Q (\values[85] [13] ), .CK (n_121_34), .D (sps__n40));
DFF_X1 \values_reg[85][14]  (.Q (\values[85] [14] ), .CK (n_121_34), .D (sps__n28));
DFF_X1 \values_reg[85][15]  (.Q (\values[85] [15] ), .CK (n_121_34), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[85]_reg  (.GCK (n_121_34), .CK (clk), .E (n_85), .SE (1'b0 ));
DFF_X1 \values_reg[86][0]  (.Q (\values[86] [0] ), .CK (n_121_33), .D (sps__n5));
DFF_X1 \values_reg[86][1]  (.Q (\values[86] [1] ), .CK (n_121_33), .D (sps__n71));
DFF_X1 \values_reg[86][2]  (.Q (\values[86] [2] ), .CK (n_121_33), .D (spc__n159));
DFF_X1 \values_reg[86][3]  (.Q (\values[86] [3] ), .CK (n_121_33), .D (sps__n78));
DFF_X1 \values_reg[86][4]  (.Q (\values[86] [4] ), .CK (n_121_33), .D (sps__n89));
DFF_X1 \values_reg[86][5]  (.Q (\values[86] [5] ), .CK (n_121_33), .D (spc__n132));
DFF_X1 \values_reg[86][6]  (.Q (\values[86] [6] ), .CK (n_121_33), .D (sps__n118));
DFF_X1 \values_reg[86][7]  (.Q (\values[86] [7] ), .CK (n_121_33), .D (spc__n127));
DFF_X1 \values_reg[86][8]  (.Q (\values[86] [8] ), .CK (n_121_33), .D (sps__n97));
DFF_X1 \values_reg[86][9]  (.Q (\values[86] [9] ), .CK (n_121_33), .D (sps__n109));
DFF_X1 \values_reg[86][10]  (.Q (\values[86] [10] ), .CK (n_121_33), .D (sps__n1));
DFF_X1 \values_reg[86][11]  (.Q (\values[86] [11] ), .CK (n_121_33), .D (sps__n12));
DFF_X1 \values_reg[86][12]  (.Q (\values[86] [12] ), .CK (n_121_33), .D (sps__n54));
DFF_X1 \values_reg[86][13]  (.Q (\values[86] [13] ), .CK (n_121_33), .D (sps__n40));
DFF_X1 \values_reg[86][14]  (.Q (\values[86] [14] ), .CK (n_121_33), .D (sps__n28));
DFF_X1 \values_reg[86][15]  (.Q (\values[86] [15] ), .CK (n_121_33), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[86]_reg  (.GCK (n_121_33), .CK (clk), .E (n_86), .SE (1'b0 ));
DFF_X1 \values_reg[87][0]  (.Q (\values[87] [0] ), .CK (n_121_32), .D (sps__n5));
DFF_X1 \values_reg[87][1]  (.Q (\values[87] [1] ), .CK (n_121_32), .D (sps__n71));
DFF_X1 \values_reg[87][2]  (.Q (\values[87] [2] ), .CK (n_121_32), .D (spc__n159));
DFF_X1 \values_reg[87][3]  (.Q (\values[87] [3] ), .CK (n_121_32), .D (sps__n78));
DFF_X1 \values_reg[87][4]  (.Q (\values[87] [4] ), .CK (n_121_32), .D (sps__n89));
DFF_X1 \values_reg[87][5]  (.Q (\values[87] [5] ), .CK (n_121_32), .D (spc__n132));
DFF_X1 \values_reg[87][6]  (.Q (\values[87] [6] ), .CK (n_121_32), .D (sps__n118));
DFF_X1 \values_reg[87][7]  (.Q (\values[87] [7] ), .CK (n_121_32), .D (spc__n127));
DFF_X1 \values_reg[87][8]  (.Q (\values[87] [8] ), .CK (n_121_32), .D (sps__n97));
DFF_X1 \values_reg[87][9]  (.Q (\values[87] [9] ), .CK (n_121_32), .D (sps__n109));
DFF_X1 \values_reg[87][10]  (.Q (\values[87] [10] ), .CK (n_121_32), .D (sps__n1));
DFF_X1 \values_reg[87][11]  (.Q (\values[87] [11] ), .CK (n_121_32), .D (sps__n12));
DFF_X1 \values_reg[87][12]  (.Q (\values[87] [12] ), .CK (n_121_32), .D (sps__n54));
DFF_X1 \values_reg[87][13]  (.Q (\values[87] [13] ), .CK (n_121_32), .D (sps__n40));
DFF_X1 \values_reg[87][14]  (.Q (\values[87] [14] ), .CK (n_121_32), .D (sps__n28));
DFF_X1 \values_reg[87][15]  (.Q (\values[87] [15] ), .CK (n_121_32), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[87]_reg  (.GCK (n_121_32), .CK (clk), .E (n_87), .SE (1'b0 ));
DFF_X1 \values_reg[88][0]  (.Q (\values[88] [0] ), .CK (n_121_31), .D (sps__n5));
DFF_X1 \values_reg[88][1]  (.Q (\values[88] [1] ), .CK (n_121_31), .D (sps__n71));
DFF_X1 \values_reg[88][2]  (.Q (\values[88] [2] ), .CK (n_121_31), .D (spc__n159));
DFF_X1 \values_reg[88][3]  (.Q (\values[88] [3] ), .CK (n_121_31), .D (sps__n77));
DFF_X1 \values_reg[88][4]  (.Q (\values[88] [4] ), .CK (n_121_31), .D (sps__n89));
DFF_X1 \values_reg[88][5]  (.Q (\values[88] [5] ), .CK (n_121_31), .D (spc__n132));
DFF_X1 \values_reg[88][6]  (.Q (\values[88] [6] ), .CK (n_121_31), .D (sps__n119));
DFF_X1 \values_reg[88][7]  (.Q (\values[88] [7] ), .CK (n_121_31), .D (spc__n127));
DFF_X1 \values_reg[88][8]  (.Q (\values[88] [8] ), .CK (n_121_31), .D (sps__n97));
DFF_X1 \values_reg[88][9]  (.Q (\values[88] [9] ), .CK (n_121_31), .D (sps__n108));
DFF_X1 \values_reg[88][10]  (.Q (\values[88] [10] ), .CK (n_121_31), .D (sps__n1));
DFF_X1 \values_reg[88][11]  (.Q (\values[88] [11] ), .CK (n_121_31), .D (sps__n11));
DFF_X1 \values_reg[88][12]  (.Q (\values[88] [12] ), .CK (n_121_31), .D (sps__n57));
DFF_X1 \values_reg[88][13]  (.Q (\values[88] [13] ), .CK (n_121_31), .D (sps__n38));
DFF_X1 \values_reg[88][14]  (.Q (\values[88] [14] ), .CK (n_121_31), .D (sps__n28));
DFF_X1 \values_reg[88][15]  (.Q (\values[88] [15] ), .CK (n_121_31), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[88]_reg  (.GCK (n_121_31), .CK (clk), .E (n_88), .SE (1'b0 ));
DFF_X1 \values_reg[89][0]  (.Q (\values[89] [0] ), .CK (n_121_30), .D (sps__n5));
DFF_X1 \values_reg[89][1]  (.Q (\values[89] [1] ), .CK (n_121_30), .D (sps__n71));
DFF_X1 \values_reg[89][2]  (.Q (\values[89] [2] ), .CK (n_121_30), .D (spc__n159));
DFF_X1 \values_reg[89][3]  (.Q (\values[89] [3] ), .CK (n_121_30), .D (sps__n77));
DFF_X1 \values_reg[89][4]  (.Q (\values[89] [4] ), .CK (n_121_30), .D (sps__n89));
DFF_X1 \values_reg[89][5]  (.Q (\values[89] [5] ), .CK (n_121_30), .D (spc__n132));
DFF_X1 \values_reg[89][6]  (.Q (\values[89] [6] ), .CK (n_121_30), .D (sps__n119));
DFF_X1 \values_reg[89][7]  (.Q (\values[89] [7] ), .CK (n_121_30), .D (spc__n127));
DFF_X1 \values_reg[89][8]  (.Q (\values[89] [8] ), .CK (n_121_30), .D (sps__n97));
DFF_X1 \values_reg[89][9]  (.Q (\values[89] [9] ), .CK (n_121_30), .D (sps__n108));
DFF_X1 \values_reg[89][10]  (.Q (\values[89] [10] ), .CK (n_121_30), .D (sps__n1));
DFF_X1 \values_reg[89][11]  (.Q (\values[89] [11] ), .CK (n_121_30), .D (sps__n11));
DFF_X1 \values_reg[89][12]  (.Q (\values[89] [12] ), .CK (n_121_30), .D (sps__n57));
DFF_X1 \values_reg[89][13]  (.Q (\values[89] [13] ), .CK (n_121_30), .D (sps__n39));
DFF_X1 \values_reg[89][14]  (.Q (\values[89] [14] ), .CK (n_121_30), .D (sps__n28));
DFF_X1 \values_reg[89][15]  (.Q (\values[89] [15] ), .CK (n_121_30), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[89]_reg  (.GCK (n_121_30), .CK (clk), .E (n_89), .SE (1'b0 ));
DFF_X1 \values_reg[90][0]  (.Q (\values[90] [0] ), .CK (n_121_29), .D (sps__n5));
DFF_X1 \values_reg[90][1]  (.Q (\values[90] [1] ), .CK (n_121_29), .D (sps__n71));
DFF_X1 \values_reg[90][2]  (.Q (\values[90] [2] ), .CK (n_121_29), .D (spc__n157));
DFF_X1 \values_reg[90][3]  (.Q (\values[90] [3] ), .CK (n_121_29), .D (sps__n79));
DFF_X1 \values_reg[90][4]  (.Q (\values[90] [4] ), .CK (n_121_29), .D (sps__n89));
DFF_X1 \values_reg[90][5]  (.Q (\values[90] [5] ), .CK (n_121_29), .D (spc__n132));
DFF_X1 \values_reg[90][6]  (.Q (\values[90] [6] ), .CK (n_121_29), .D (sps__n118));
DFF_X1 \values_reg[90][7]  (.Q (\values[90] [7] ), .CK (n_121_29), .D (spc__n126));
DFF_X1 \values_reg[90][8]  (.Q (\values[90] [8] ), .CK (n_121_29), .D (sps__n97));
DFF_X1 \values_reg[90][9]  (.Q (\values[90] [9] ), .CK (n_121_29), .D (sps__n109));
DFF_X1 \values_reg[90][10]  (.Q (\values[90] [10] ), .CK (n_121_29), .D (sps__n1));
DFF_X1 \values_reg[90][11]  (.Q (\values[90] [11] ), .CK (n_121_29), .D (sps__n12));
DFF_X1 \values_reg[90][12]  (.Q (\values[90] [12] ), .CK (n_121_29), .D (sps__n55));
DFF_X1 \values_reg[90][13]  (.Q (\values[90] [13] ), .CK (n_121_29), .D (sps__n40));
DFF_X1 \values_reg[90][14]  (.Q (\values[90] [14] ), .CK (n_121_29), .D (sps__n28));
DFF_X1 \values_reg[90][15]  (.Q (\values[90] [15] ), .CK (n_121_29), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[90]_reg  (.GCK (n_121_29), .CK (clk), .E (n_90), .SE (1'b0 ));
DFF_X1 \values_reg[91][0]  (.Q (\values[91] [0] ), .CK (n_121_28), .D (sps__n5));
DFF_X1 \values_reg[91][1]  (.Q (\values[91] [1] ), .CK (n_121_28), .D (sps__n71));
DFF_X1 \values_reg[91][2]  (.Q (\values[91] [2] ), .CK (n_121_28), .D (spc__n157));
DFF_X1 \values_reg[91][3]  (.Q (\values[91] [3] ), .CK (n_121_28), .D (sps__n79));
DFF_X1 \values_reg[91][4]  (.Q (\values[91] [4] ), .CK (n_121_28), .D (sps__n89));
DFF_X1 \values_reg[91][5]  (.Q (\values[91] [5] ), .CK (n_121_28), .D (spc__n132));
DFF_X1 \values_reg[91][6]  (.Q (\values[91] [6] ), .CK (n_121_28), .D (sps__n118));
DFF_X1 \values_reg[91][7]  (.Q (\values[91] [7] ), .CK (n_121_28), .D (spc__n126));
DFF_X1 \values_reg[91][8]  (.Q (\values[91] [8] ), .CK (n_121_28), .D (sps__n97));
DFF_X1 \values_reg[91][9]  (.Q (\values[91] [9] ), .CK (n_121_28), .D (sps__n109));
DFF_X1 \values_reg[91][10]  (.Q (\values[91] [10] ), .CK (n_121_28), .D (sps__n1));
DFF_X1 \values_reg[91][11]  (.Q (\values[91] [11] ), .CK (n_121_28), .D (sps__n12));
DFF_X1 \values_reg[91][12]  (.Q (\values[91] [12] ), .CK (n_121_28), .D (sps__n55));
DFF_X1 \values_reg[91][13]  (.Q (\values[91] [13] ), .CK (n_121_28), .D (sps__n40));
DFF_X1 \values_reg[91][14]  (.Q (\values[91] [14] ), .CK (n_121_28), .D (sps__n28));
DFF_X1 \values_reg[91][15]  (.Q (\values[91] [15] ), .CK (n_121_28), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[91]_reg  (.GCK (n_121_28), .CK (clk), .E (n_91), .SE (1'b0 ));
DFF_X1 \values_reg[92][0]  (.Q (\values[92] [0] ), .CK (n_121_27), .D (sps__n5));
DFF_X1 \values_reg[92][1]  (.Q (\values[92] [1] ), .CK (n_121_27), .D (sps__n71));
DFF_X1 \values_reg[92][2]  (.Q (\values[92] [2] ), .CK (n_121_27), .D (spc__n159));
DFF_X1 \values_reg[92][3]  (.Q (\values[92] [3] ), .CK (n_121_27), .D (sps__n77));
DFF_X1 \values_reg[92][4]  (.Q (\values[92] [4] ), .CK (n_121_27), .D (sps__n89));
DFF_X1 \values_reg[92][5]  (.Q (\values[92] [5] ), .CK (n_121_27), .D (spc__n132));
DFF_X1 \values_reg[92][6]  (.Q (\values[92] [6] ), .CK (n_121_27), .D (sps__n119));
DFF_X1 \values_reg[92][7]  (.Q (\values[92] [7] ), .CK (n_121_27), .D (spc__n127));
DFF_X1 \values_reg[92][8]  (.Q (\values[92] [8] ), .CK (n_121_27), .D (sps__n97));
DFF_X1 \values_reg[92][9]  (.Q (\values[92] [9] ), .CK (n_121_27), .D (sps__n108));
DFF_X1 \values_reg[92][10]  (.Q (\values[92] [10] ), .CK (n_121_27), .D (sps__n1));
DFF_X1 \values_reg[92][11]  (.Q (\values[92] [11] ), .CK (n_121_27), .D (sps__n12));
DFF_X1 \values_reg[92][12]  (.Q (\values[92] [12] ), .CK (n_121_27), .D (sps__n57));
DFF_X1 \values_reg[92][13]  (.Q (\values[92] [13] ), .CK (n_121_27), .D (sps__n39));
DFF_X1 \values_reg[92][14]  (.Q (\values[92] [14] ), .CK (n_121_27), .D (sps__n28));
DFF_X1 \values_reg[92][15]  (.Q (\values[92] [15] ), .CK (n_121_27), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[92]_reg  (.GCK (n_121_27), .CK (clk), .E (n_92), .SE (1'b0 ));
DFF_X1 \values_reg[93][0]  (.Q (\values[93] [0] ), .CK (n_121_26), .D (sps__n5));
DFF_X1 \values_reg[93][1]  (.Q (\values[93] [1] ), .CK (n_121_26), .D (sps__n71));
DFF_X1 \values_reg[93][2]  (.Q (\values[93] [2] ), .CK (n_121_26), .D (spc__n159));
DFF_X1 \values_reg[93][3]  (.Q (\values[93] [3] ), .CK (n_121_26), .D (sps__n78));
DFF_X1 \values_reg[93][4]  (.Q (\values[93] [4] ), .CK (n_121_26), .D (sps__n89));
DFF_X1 \values_reg[93][5]  (.Q (\values[93] [5] ), .CK (n_121_26), .D (spc__n132));
DFF_X1 \values_reg[93][6]  (.Q (\values[93] [6] ), .CK (n_121_26), .D (sps__n118));
DFF_X1 \values_reg[93][7]  (.Q (\values[93] [7] ), .CK (n_121_26), .D (spc__n127));
DFF_X1 \values_reg[93][8]  (.Q (\values[93] [8] ), .CK (n_121_26), .D (sps__n97));
DFF_X1 \values_reg[93][9]  (.Q (\values[93] [9] ), .CK (n_121_26), .D (sps__n109));
DFF_X1 \values_reg[93][10]  (.Q (\values[93] [10] ), .CK (n_121_26), .D (sps__n1));
DFF_X1 \values_reg[93][11]  (.Q (\values[93] [11] ), .CK (n_121_26), .D (sps__n12));
DFF_X1 \values_reg[93][12]  (.Q (\values[93] [12] ), .CK (n_121_26), .D (sps__n54));
DFF_X1 \values_reg[93][13]  (.Q (\values[93] [13] ), .CK (n_121_26), .D (sps__n40));
DFF_X1 \values_reg[93][14]  (.Q (\values[93] [14] ), .CK (n_121_26), .D (sps__n28));
DFF_X1 \values_reg[93][15]  (.Q (\values[93] [15] ), .CK (n_121_26), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[93]_reg  (.GCK (n_121_26), .CK (clk), .E (n_93), .SE (1'b0 ));
DFF_X1 \values_reg[94][0]  (.Q (\values[94] [0] ), .CK (n_121_25), .D (sps__n5));
DFF_X1 \values_reg[94][1]  (.Q (\values[94] [1] ), .CK (n_121_25), .D (sps__n71));
DFF_X1 \values_reg[94][2]  (.Q (\values[94] [2] ), .CK (n_121_25), .D (spc__n157));
DFF_X1 \values_reg[94][3]  (.Q (\values[94] [3] ), .CK (n_121_25), .D (sps__n79));
DFF_X1 \values_reg[94][4]  (.Q (\values[94] [4] ), .CK (n_121_25), .D (sps__n89));
DFF_X1 \values_reg[94][5]  (.Q (\values[94] [5] ), .CK (n_121_25), .D (spc__n132));
DFF_X1 \values_reg[94][6]  (.Q (\values[94] [6] ), .CK (n_121_25), .D (sps__n118));
DFF_X1 \values_reg[94][7]  (.Q (\values[94] [7] ), .CK (n_121_25), .D (spc__n126));
DFF_X1 \values_reg[94][8]  (.Q (\values[94] [8] ), .CK (n_121_25), .D (sps__n97));
DFF_X1 \values_reg[94][9]  (.Q (\values[94] [9] ), .CK (n_121_25), .D (sps__n109));
DFF_X1 \values_reg[94][10]  (.Q (\values[94] [10] ), .CK (n_121_25), .D (sps__n1));
DFF_X1 \values_reg[94][11]  (.Q (\values[94] [11] ), .CK (n_121_25), .D (sps__n12));
DFF_X1 \values_reg[94][12]  (.Q (\values[94] [12] ), .CK (n_121_25), .D (sps__n55));
DFF_X1 \values_reg[94][13]  (.Q (\values[94] [13] ), .CK (n_121_25), .D (sps__n40));
DFF_X1 \values_reg[94][14]  (.Q (\values[94] [14] ), .CK (n_121_25), .D (sps__n28));
DFF_X1 \values_reg[94][15]  (.Q (\values[94] [15] ), .CK (n_121_25), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[94]_reg  (.GCK (n_121_25), .CK (clk), .E (n_94), .SE (1'b0 ));
DFF_X1 \values_reg[95][0]  (.Q (\values[95] [0] ), .CK (n_121_24), .D (sps__n5));
DFF_X1 \values_reg[95][1]  (.Q (\values[95] [1] ), .CK (n_121_24), .D (sps__n71));
DFF_X1 \values_reg[95][2]  (.Q (\values[95] [2] ), .CK (n_121_24), .D (spc__n157));
DFF_X1 \values_reg[95][3]  (.Q (\values[95] [3] ), .CK (n_121_24), .D (sps__n79));
DFF_X1 \values_reg[95][4]  (.Q (\values[95] [4] ), .CK (n_121_24), .D (sps__n89));
DFF_X1 \values_reg[95][5]  (.Q (\values[95] [5] ), .CK (n_121_24), .D (spc__n132));
DFF_X1 \values_reg[95][6]  (.Q (\values[95] [6] ), .CK (n_121_24), .D (sps__n118));
DFF_X1 \values_reg[95][7]  (.Q (\values[95] [7] ), .CK (n_121_24), .D (spc__n126));
DFF_X1 \values_reg[95][8]  (.Q (\values[95] [8] ), .CK (n_121_24), .D (sps__n97));
DFF_X1 \values_reg[95][9]  (.Q (\values[95] [9] ), .CK (n_121_24), .D (sps__n109));
DFF_X1 \values_reg[95][10]  (.Q (\values[95] [10] ), .CK (n_121_24), .D (sps__n1));
DFF_X1 \values_reg[95][11]  (.Q (\values[95] [11] ), .CK (n_121_24), .D (sps__n12));
DFF_X1 \values_reg[95][12]  (.Q (\values[95] [12] ), .CK (n_121_24), .D (sps__n55));
DFF_X1 \values_reg[95][13]  (.Q (\values[95] [13] ), .CK (n_121_24), .D (sps__n40));
DFF_X1 \values_reg[95][14]  (.Q (\values[95] [14] ), .CK (n_121_24), .D (sps__n28));
DFF_X1 \values_reg[95][15]  (.Q (\values[95] [15] ), .CK (n_121_24), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[95]_reg  (.GCK (n_121_24), .CK (clk), .E (n_95), .SE (1'b0 ));
DFF_X1 \values_reg[96][0]  (.Q (\values[96] [0] ), .CK (n_121_23), .D (sps__n5));
DFF_X1 \values_reg[96][1]  (.Q (\values[96] [1] ), .CK (n_121_23), .D (sps__n71));
DFF_X1 \values_reg[96][2]  (.Q (\values[96] [2] ), .CK (n_121_23), .D (spc__n157));
DFF_X1 \values_reg[96][3]  (.Q (\values[96] [3] ), .CK (n_121_23), .D (sps__n79));
DFF_X1 \values_reg[96][4]  (.Q (\values[96] [4] ), .CK (n_121_23), .D (sps__n89));
DFF_X1 \values_reg[96][5]  (.Q (\values[96] [5] ), .CK (n_121_23), .D (spc__n132));
DFF_X1 \values_reg[96][6]  (.Q (\values[96] [6] ), .CK (n_121_23), .D (sps__n118));
DFF_X1 \values_reg[96][7]  (.Q (\values[96] [7] ), .CK (n_121_23), .D (spc__n126));
DFF_X1 \values_reg[96][8]  (.Q (\values[96] [8] ), .CK (n_121_23), .D (sps__n97));
DFF_X1 \values_reg[96][9]  (.Q (\values[96] [9] ), .CK (n_121_23), .D (sps__n109));
DFF_X1 \values_reg[96][10]  (.Q (\values[96] [10] ), .CK (n_121_23), .D (sps__n1));
DFF_X1 \values_reg[96][11]  (.Q (\values[96] [11] ), .CK (n_121_23), .D (sps__n12));
DFF_X1 \values_reg[96][12]  (.Q (\values[96] [12] ), .CK (n_121_23), .D (sps__n55));
DFF_X1 \values_reg[96][13]  (.Q (\values[96] [13] ), .CK (n_121_23), .D (sps__n40));
DFF_X1 \values_reg[96][14]  (.Q (\values[96] [14] ), .CK (n_121_23), .D (sps__n28));
DFF_X1 \values_reg[96][15]  (.Q (\values[96] [15] ), .CK (n_121_23), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[96]_reg  (.GCK (n_121_23), .CK (clk), .E (n_96), .SE (1'b0 ));
DFF_X1 \values_reg[25][0]  (.Q (\values[25] [0] ), .CK (n_121_22), .D (sps__n5));
DFF_X1 \values_reg[25][1]  (.Q (\values[25] [1] ), .CK (n_121_22), .D (sps__n71));
DFF_X1 \values_reg[25][2]  (.Q (\values[25] [2] ), .CK (n_121_22), .D (spc__n159));
DFF_X1 \values_reg[25][3]  (.Q (\values[25] [3] ), .CK (n_121_22), .D (sps__n77));
DFF_X1 \values_reg[25][4]  (.Q (\values[25] [4] ), .CK (n_121_22), .D (sps__n89));
DFF_X1 \values_reg[25][5]  (.Q (\values[25] [5] ), .CK (n_121_22), .D (spc__n132));
DFF_X1 \values_reg[25][6]  (.Q (\values[25] [6] ), .CK (n_121_22), .D (sps__n117));
DFF_X1 \values_reg[25][7]  (.Q (\values[25] [7] ), .CK (n_121_22), .D (spc__n127));
DFF_X1 \values_reg[25][8]  (.Q (\values[25] [8] ), .CK (n_121_22), .D (sps__n97));
DFF_X1 \values_reg[25][9]  (.Q (\values[25] [9] ), .CK (n_121_22), .D (sps__n108));
DFF_X1 \values_reg[25][10]  (.Q (\values[25] [10] ), .CK (n_121_22), .D (sps__n1));
DFF_X1 \values_reg[25][11]  (.Q (\values[25] [11] ), .CK (n_121_22), .D (sps__n12));
DFF_X1 \values_reg[25][12]  (.Q (\values[25] [12] ), .CK (n_121_22), .D (sps__n57));
DFF_X1 \values_reg[25][13]  (.Q (\values[25] [13] ), .CK (n_121_22), .D (sps__n39));
DFF_X1 \values_reg[25][14]  (.Q (\values[25] [14] ), .CK (n_121_22), .D (sps__n25));
DFF_X1 \values_reg[25][15]  (.Q (\values[25] [15] ), .CK (n_121_22), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[25]_reg  (.GCK (n_121_22), .CK (clk), .E (n_25), .SE (1'b0 ));
DFF_X1 \values_reg[24][0]  (.Q (\values[24] [0] ), .CK (n_121_21), .D (sps__n5));
DFF_X1 \values_reg[24][1]  (.Q (\values[24] [1] ), .CK (n_121_21), .D (sps__n71));
DFF_X1 \values_reg[24][2]  (.Q (\values[24] [2] ), .CK (n_121_21), .D (spc__n159));
DFF_X1 \values_reg[24][3]  (.Q (\values[24] [3] ), .CK (n_121_21), .D (sps__n77));
DFF_X1 \values_reg[24][4]  (.Q (\values[24] [4] ), .CK (n_121_21), .D (sps__n90));
DFF_X1 \values_reg[24][5]  (.Q (\values[24] [5] ), .CK (n_121_21), .D (spc__n132));
DFF_X1 \values_reg[24][6]  (.Q (\values[24] [6] ), .CK (n_121_21), .D (sps__n117));
DFF_X1 \values_reg[24][7]  (.Q (\values[24] [7] ), .CK (n_121_21), .D (spc__n127));
DFF_X1 \values_reg[24][8]  (.Q (\values[24] [8] ), .CK (n_121_21), .D (sps__n97));
DFF_X1 \values_reg[24][9]  (.Q (\values[24] [9] ), .CK (n_121_21), .D (sps__n108));
DFF_X1 \values_reg[24][10]  (.Q (\values[24] [10] ), .CK (n_121_21), .D (sps__n1));
DFF_X1 \values_reg[24][11]  (.Q (\values[24] [11] ), .CK (n_121_21), .D (sps__n12));
DFF_X1 \values_reg[24][12]  (.Q (\values[24] [12] ), .CK (n_121_21), .D (sps__n57));
DFF_X1 \values_reg[24][13]  (.Q (\values[24] [13] ), .CK (n_121_21), .D (sps__n40));
DFF_X1 \values_reg[24][14]  (.Q (\values[24] [14] ), .CK (n_121_21), .D (sps__n25));
DFF_X1 \values_reg[24][15]  (.Q (\values[24] [15] ), .CK (n_121_21), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[24]_reg  (.GCK (n_121_21), .CK (clk), .E (n_24), .SE (1'b0 ));
DFF_X1 \values_reg[23][0]  (.Q (\values[23] [0] ), .CK (n_121_20), .D (sps__n5));
DFF_X1 \values_reg[23][1]  (.Q (\values[23] [1] ), .CK (n_121_20), .D (sps__n71));
DFF_X1 \values_reg[23][2]  (.Q (\values[23] [2] ), .CK (n_121_20), .D (spc__n159));
DFF_X1 \values_reg[23][3]  (.Q (\values[23] [3] ), .CK (n_121_20), .D (sps__n78));
DFF_X1 \values_reg[23][4]  (.Q (\values[23] [4] ), .CK (n_121_20), .D (sps__n89));
DFF_X1 \values_reg[23][5]  (.Q (\values[23] [5] ), .CK (n_121_20), .D (spc__n132));
DFF_X1 \values_reg[23][6]  (.Q (\values[23] [6] ), .CK (n_121_20), .D (sps__n118));
DFF_X1 \values_reg[23][7]  (.Q (\values[23] [7] ), .CK (n_121_20), .D (spc__n127));
DFF_X1 \values_reg[23][8]  (.Q (\values[23] [8] ), .CK (n_121_20), .D (sps__n97));
DFF_X1 \values_reg[23][9]  (.Q (\values[23] [9] ), .CK (n_121_20), .D (sps__n109));
DFF_X1 \values_reg[23][10]  (.Q (\values[23] [10] ), .CK (n_121_20), .D (sps__n1));
DFF_X1 \values_reg[23][11]  (.Q (\values[23] [11] ), .CK (n_121_20), .D (sps__n12));
DFF_X1 \values_reg[23][12]  (.Q (\values[23] [12] ), .CK (n_121_20), .D (sps__n54));
DFF_X1 \values_reg[23][13]  (.Q (\values[23] [13] ), .CK (n_121_20), .D (sps__n40));
DFF_X1 \values_reg[23][14]  (.Q (\values[23] [14] ), .CK (n_121_20), .D (sps__n28));
DFF_X1 \values_reg[23][15]  (.Q (\values[23] [15] ), .CK (n_121_20), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[23]_reg  (.GCK (n_121_20), .CK (clk), .E (n_23), .SE (1'b0 ));
DFF_X1 \values_reg[22][0]  (.Q (\values[22] [0] ), .CK (n_121_19), .D (sps__n5));
DFF_X1 \values_reg[22][1]  (.Q (\values[22] [1] ), .CK (n_121_19), .D (sps__n71));
DFF_X1 \values_reg[22][2]  (.Q (\values[22] [2] ), .CK (n_121_19), .D (spc__n159));
DFF_X1 \values_reg[22][3]  (.Q (\values[22] [3] ), .CK (n_121_19), .D (sps__n77));
DFF_X1 \values_reg[22][4]  (.Q (\values[22] [4] ), .CK (n_121_19), .D (sps__n89));
DFF_X1 \values_reg[22][5]  (.Q (\values[22] [5] ), .CK (n_121_19), .D (spc__n132));
DFF_X1 \values_reg[22][6]  (.Q (\values[22] [6] ), .CK (n_121_19), .D (sps__n117));
DFF_X1 \values_reg[22][7]  (.Q (\values[22] [7] ), .CK (n_121_19), .D (spc__n127));
DFF_X1 \values_reg[22][8]  (.Q (\values[22] [8] ), .CK (n_121_19), .D (sps__n97));
DFF_X1 \values_reg[22][9]  (.Q (\values[22] [9] ), .CK (n_121_19), .D (sps__n109));
DFF_X1 \values_reg[22][10]  (.Q (\values[22] [10] ), .CK (n_121_19), .D (sps__n1));
DFF_X1 \values_reg[22][11]  (.Q (\values[22] [11] ), .CK (n_121_19), .D (sps__n12));
DFF_X1 \values_reg[22][12]  (.Q (\values[22] [12] ), .CK (n_121_19), .D (sps__n54));
DFF_X1 \values_reg[22][13]  (.Q (\values[22] [13] ), .CK (n_121_19), .D (sps__n39));
DFF_X1 \values_reg[22][14]  (.Q (\values[22] [14] ), .CK (n_121_19), .D (sps__n27));
DFF_X1 \values_reg[22][15]  (.Q (\values[22] [15] ), .CK (n_121_19), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[22]_reg  (.GCK (n_121_19), .CK (clk), .E (n_22), .SE (1'b0 ));
DFF_X1 \values_reg[21][0]  (.Q (\values[21] [0] ), .CK (n_121_18), .D (sps__n5));
DFF_X1 \values_reg[21][1]  (.Q (\values[21] [1] ), .CK (n_121_18), .D (sps__n71));
DFF_X1 \values_reg[21][2]  (.Q (\values[21] [2] ), .CK (n_121_18), .D (spc__n159));
DFF_X1 \values_reg[21][3]  (.Q (\values[21] [3] ), .CK (n_121_18), .D (sps__n77));
DFF_X1 \values_reg[21][4]  (.Q (\values[21] [4] ), .CK (n_121_18), .D (sps__n89));
DFF_X1 \values_reg[21][5]  (.Q (\values[21] [5] ), .CK (n_121_18), .D (spc__n132));
DFF_X1 \values_reg[21][6]  (.Q (\values[21] [6] ), .CK (n_121_18), .D (sps__n118));
DFF_X1 \values_reg[21][7]  (.Q (\values[21] [7] ), .CK (n_121_18), .D (spc__n127));
DFF_X1 \values_reg[21][8]  (.Q (\values[21] [8] ), .CK (n_121_18), .D (sps__n97));
DFF_X1 \values_reg[21][9]  (.Q (\values[21] [9] ), .CK (n_121_18), .D (sps__n109));
DFF_X1 \values_reg[21][10]  (.Q (\values[21] [10] ), .CK (n_121_18), .D (sps__n1));
DFF_X1 \values_reg[21][11]  (.Q (\values[21] [11] ), .CK (n_121_18), .D (sps__n12));
DFF_X1 \values_reg[21][12]  (.Q (\values[21] [12] ), .CK (n_121_18), .D (sps__n54));
DFF_X1 \values_reg[21][13]  (.Q (\values[21] [13] ), .CK (n_121_18), .D (sps__n39));
DFF_X1 \values_reg[21][14]  (.Q (\values[21] [14] ), .CK (n_121_18), .D (sps__n27));
DFF_X1 \values_reg[21][15]  (.Q (\values[21] [15] ), .CK (n_121_18), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[21]_reg  (.GCK (n_121_18), .CK (clk), .E (n_21), .SE (1'b0 ));
DFF_X1 \values_reg[20][0]  (.Q (\values[20] [0] ), .CK (n_121_17), .D (sps__n5));
DFF_X1 \values_reg[20][1]  (.Q (\values[20] [1] ), .CK (n_121_17), .D (sps__n71));
DFF_X1 \values_reg[20][2]  (.Q (\values[20] [2] ), .CK (n_121_17), .D (spc__n159));
DFF_X1 \values_reg[20][3]  (.Q (\values[20] [3] ), .CK (n_121_17), .D (sps__n77));
DFF_X1 \values_reg[20][4]  (.Q (\values[20] [4] ), .CK (n_121_17), .D (sps__n89));
DFF_X1 \values_reg[20][5]  (.Q (\values[20] [5] ), .CK (n_121_17), .D (spc__n132));
DFF_X1 \values_reg[20][6]  (.Q (\values[20] [6] ), .CK (n_121_17), .D (sps__n117));
DFF_X1 \values_reg[20][7]  (.Q (\values[20] [7] ), .CK (n_121_17), .D (spc__n127));
DFF_X1 \values_reg[20][8]  (.Q (\values[20] [8] ), .CK (n_121_17), .D (sps__n97));
DFF_X1 \values_reg[20][9]  (.Q (\values[20] [9] ), .CK (n_121_17), .D (sps__n108));
DFF_X1 \values_reg[20][10]  (.Q (\values[20] [10] ), .CK (n_121_17), .D (sps__n1));
DFF_X1 \values_reg[20][11]  (.Q (\values[20] [11] ), .CK (n_121_17), .D (sps__n12));
DFF_X1 \values_reg[20][12]  (.Q (\values[20] [12] ), .CK (n_121_17), .D (sps__n57));
DFF_X1 \values_reg[20][13]  (.Q (\values[20] [13] ), .CK (n_121_17), .D (sps__n40));
DFF_X1 \values_reg[20][14]  (.Q (\values[20] [14] ), .CK (n_121_17), .D (sps__n25));
DFF_X1 \values_reg[20][15]  (.Q (\values[20] [15] ), .CK (n_121_17), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[20]_reg  (.GCK (n_121_17), .CK (clk), .E (n_20), .SE (1'b0 ));
DFF_X1 \values_reg[19][0]  (.Q (\values[19] [0] ), .CK (n_121_16), .D (sps__n5));
DFF_X1 \values_reg[19][1]  (.Q (\values[19] [1] ), .CK (n_121_16), .D (sps__n71));
DFF_X1 \values_reg[19][2]  (.Q (\values[19] [2] ), .CK (n_121_16), .D (spc__n159));
DFF_X1 \values_reg[19][3]  (.Q (\values[19] [3] ), .CK (n_121_16), .D (sps__n77));
DFF_X1 \values_reg[19][4]  (.Q (\values[19] [4] ), .CK (n_121_16), .D (sps__n89));
DFF_X1 \values_reg[19][5]  (.Q (\values[19] [5] ), .CK (n_121_16), .D (spc__n132));
DFF_X1 \values_reg[19][6]  (.Q (\values[19] [6] ), .CK (n_121_16), .D (sps__n118));
DFF_X1 \values_reg[19][7]  (.Q (\values[19] [7] ), .CK (n_121_16), .D (spc__n127));
DFF_X1 \values_reg[19][8]  (.Q (\values[19] [8] ), .CK (n_121_16), .D (sps__n97));
DFF_X1 \values_reg[19][9]  (.Q (\values[19] [9] ), .CK (n_121_16), .D (sps__n109));
DFF_X1 \values_reg[19][10]  (.Q (\values[19] [10] ), .CK (n_121_16), .D (sps__n1));
DFF_X1 \values_reg[19][11]  (.Q (\values[19] [11] ), .CK (n_121_16), .D (sps__n12));
DFF_X1 \values_reg[19][12]  (.Q (\values[19] [12] ), .CK (n_121_16), .D (sps__n54));
DFF_X1 \values_reg[19][13]  (.Q (\values[19] [13] ), .CK (n_121_16), .D (sps__n40));
DFF_X1 \values_reg[19][14]  (.Q (\values[19] [14] ), .CK (n_121_16), .D (sps__n27));
DFF_X1 \values_reg[19][15]  (.Q (\values[19] [15] ), .CK (n_121_16), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[19]_reg  (.GCK (n_121_16), .CK (clk), .E (n_19), .SE (1'b0 ));
DFF_X1 \values_reg[18][0]  (.Q (\values[18] [0] ), .CK (n_121_15), .D (sps__n5));
DFF_X1 \values_reg[18][1]  (.Q (\values[18] [1] ), .CK (n_121_15), .D (sps__n71));
DFF_X1 \values_reg[18][2]  (.Q (\values[18] [2] ), .CK (n_121_15), .D (spc__n159));
DFF_X1 \values_reg[18][3]  (.Q (\values[18] [3] ), .CK (n_121_15), .D (sps__n77));
DFF_X1 \values_reg[18][4]  (.Q (\values[18] [4] ), .CK (n_121_15), .D (sps__n89));
DFF_X1 \values_reg[18][5]  (.Q (\values[18] [5] ), .CK (n_121_15), .D (spc__n132));
DFF_X1 \values_reg[18][6]  (.Q (\values[18] [6] ), .CK (n_121_15), .D (sps__n118));
DFF_X1 \values_reg[18][7]  (.Q (\values[18] [7] ), .CK (n_121_15), .D (spc__n127));
DFF_X1 \values_reg[18][8]  (.Q (\values[18] [8] ), .CK (n_121_15), .D (sps__n97));
DFF_X1 \values_reg[18][9]  (.Q (\values[18] [9] ), .CK (n_121_15), .D (sps__n109));
DFF_X1 \values_reg[18][10]  (.Q (\values[18] [10] ), .CK (n_121_15), .D (sps__n1));
DFF_X1 \values_reg[18][11]  (.Q (\values[18] [11] ), .CK (n_121_15), .D (sps__n12));
DFF_X1 \values_reg[18][12]  (.Q (\values[18] [12] ), .CK (n_121_15), .D (sps__n54));
DFF_X1 \values_reg[18][13]  (.Q (\values[18] [13] ), .CK (n_121_15), .D (sps__n39));
DFF_X1 \values_reg[18][14]  (.Q (\values[18] [14] ), .CK (n_121_15), .D (sps__n27));
DFF_X1 \values_reg[18][15]  (.Q (\values[18] [15] ), .CK (n_121_15), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[18]_reg  (.GCK (n_121_15), .CK (clk), .E (n_18), .SE (1'b0 ));
DFF_X1 \values_reg[17][0]  (.Q (\values[17] [0] ), .CK (n_121_14), .D (sps__n5));
DFF_X1 \values_reg[17][1]  (.Q (\values[17] [1] ), .CK (n_121_14), .D (sps__n71));
DFF_X1 \values_reg[17][2]  (.Q (\values[17] [2] ), .CK (n_121_14), .D (spc__n159));
DFF_X1 \values_reg[17][3]  (.Q (\values[17] [3] ), .CK (n_121_14), .D (sps__n77));
DFF_X1 \values_reg[17][4]  (.Q (\values[17] [4] ), .CK (n_121_14), .D (sps__n89));
DFF_X1 \values_reg[17][5]  (.Q (\values[17] [5] ), .CK (n_121_14), .D (spc__n132));
DFF_X1 \values_reg[17][6]  (.Q (\values[17] [6] ), .CK (n_121_14), .D (sps__n117));
DFF_X1 \values_reg[17][7]  (.Q (\values[17] [7] ), .CK (n_121_14), .D (spc__n127));
DFF_X1 \values_reg[17][8]  (.Q (\values[17] [8] ), .CK (n_121_14), .D (sps__n97));
DFF_X1 \values_reg[17][9]  (.Q (\values[17] [9] ), .CK (n_121_14), .D (sps__n108));
DFF_X1 \values_reg[17][10]  (.Q (\values[17] [10] ), .CK (n_121_14), .D (sps__n1));
DFF_X1 \values_reg[17][11]  (.Q (\values[17] [11] ), .CK (n_121_14), .D (sps__n10));
DFF_X1 \values_reg[17][12]  (.Q (\values[17] [12] ), .CK (n_121_14), .D (sps__n54));
DFF_X1 \values_reg[17][13]  (.Q (\values[17] [13] ), .CK (n_121_14), .D (sps__n39));
DFF_X1 \values_reg[17][14]  (.Q (\values[17] [14] ), .CK (n_121_14), .D (sps__n27));
DFF_X1 \values_reg[17][15]  (.Q (\values[17] [15] ), .CK (n_121_14), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[17]_reg  (.GCK (n_121_14), .CK (clk), .E (n_17), .SE (1'b0 ));
DFF_X1 \values_reg[16][0]  (.Q (\values[16] [0] ), .CK (n_121_13), .D (sps__n5));
DFF_X1 \values_reg[16][1]  (.Q (\values[16] [1] ), .CK (n_121_13), .D (sps__n71));
DFF_X1 \values_reg[16][2]  (.Q (\values[16] [2] ), .CK (n_121_13), .D (spc__n159));
DFF_X1 \values_reg[16][3]  (.Q (\values[16] [3] ), .CK (n_121_13), .D (sps__n77));
DFF_X1 \values_reg[16][4]  (.Q (\values[16] [4] ), .CK (n_121_13), .D (sps__n90));
DFF_X1 \values_reg[16][5]  (.Q (\values[16] [5] ), .CK (n_121_13), .D (spc__n132));
DFF_X1 \values_reg[16][6]  (.Q (\values[16] [6] ), .CK (n_121_13), .D (sps__n117));
DFF_X1 \values_reg[16][7]  (.Q (\values[16] [7] ), .CK (n_121_13), .D (spc__n127));
DFF_X1 \values_reg[16][8]  (.Q (\values[16] [8] ), .CK (n_121_13), .D (sps__n97));
DFF_X1 \values_reg[16][9]  (.Q (\values[16] [9] ), .CK (n_121_13), .D (sps__n108));
DFF_X1 \values_reg[16][10]  (.Q (\values[16] [10] ), .CK (n_121_13), .D (sps__n1));
DFF_X1 \values_reg[16][11]  (.Q (\values[16] [11] ), .CK (n_121_13), .D (sps__n12));
DFF_X1 \values_reg[16][12]  (.Q (\values[16] [12] ), .CK (n_121_13), .D (sps__n54));
DFF_X1 \values_reg[16][13]  (.Q (\values[16] [13] ), .CK (n_121_13), .D (sps__n39));
DFF_X1 \values_reg[16][14]  (.Q (\values[16] [14] ), .CK (n_121_13), .D (sps__n27));
DFF_X1 \values_reg[16][15]  (.Q (\values[16] [15] ), .CK (n_121_13), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[16]_reg  (.GCK (n_121_13), .CK (clk), .E (n_16), .SE (1'b0 ));
DFF_X1 \values_reg[15][0]  (.Q (\values[15] [0] ), .CK (n_121_12), .D (sps__n5));
DFF_X1 \values_reg[15][1]  (.Q (\values[15] [1] ), .CK (n_121_12), .D (sps__n71));
DFF_X1 \values_reg[15][2]  (.Q (\values[15] [2] ), .CK (n_121_12), .D (spc__n159));
DFF_X1 \values_reg[15][3]  (.Q (\values[15] [3] ), .CK (n_121_12), .D (sps__n77));
DFF_X1 \values_reg[15][4]  (.Q (\values[15] [4] ), .CK (n_121_12), .D (sps__n90));
DFF_X1 \values_reg[15][5]  (.Q (\values[15] [5] ), .CK (n_121_12), .D (spc__n132));
DFF_X1 \values_reg[15][6]  (.Q (\values[15] [6] ), .CK (n_121_12), .D (sps__n117));
DFF_X1 \values_reg[15][7]  (.Q (\values[15] [7] ), .CK (n_121_12), .D (spc__n127));
DFF_X1 \values_reg[15][8]  (.Q (\values[15] [8] ), .CK (n_121_12), .D (sps__n97));
DFF_X1 \values_reg[15][9]  (.Q (\values[15] [9] ), .CK (n_121_12), .D (sps__n110));
DFF_X1 \values_reg[15][10]  (.Q (\values[15] [10] ), .CK (n_121_12), .D (sps__n1));
DFF_X1 \values_reg[15][11]  (.Q (\values[15] [11] ), .CK (n_121_12), .D (sps__n11));
DFF_X1 \values_reg[15][12]  (.Q (\values[15] [12] ), .CK (n_121_12), .D (sps__n57));
DFF_X1 \values_reg[15][13]  (.Q (\values[15] [13] ), .CK (n_121_12), .D (sps__n38));
DFF_X1 \values_reg[15][14]  (.Q (\values[15] [14] ), .CK (n_121_12), .D (sps__n28));
DFF_X1 \values_reg[15][15]  (.Q (\values[15] [15] ), .CK (n_121_12), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[15]_reg  (.GCK (n_121_12), .CK (clk), .E (n_15), .SE (1'b0 ));
DFF_X1 \values_reg[14][0]  (.Q (\values[14] [0] ), .CK (n_121_11), .D (sps__n5));
DFF_X1 \values_reg[14][1]  (.Q (\values[14] [1] ), .CK (n_121_11), .D (sps__n71));
DFF_X1 \values_reg[14][2]  (.Q (\values[14] [2] ), .CK (n_121_11), .D (spc__n159));
DFF_X1 \values_reg[14][3]  (.Q (\values[14] [3] ), .CK (n_121_11), .D (sps__n77));
DFF_X1 \values_reg[14][4]  (.Q (\values[14] [4] ), .CK (n_121_11), .D (sps__n90));
DFF_X1 \values_reg[14][5]  (.Q (\values[14] [5] ), .CK (n_121_11), .D (spc__n132));
DFF_X1 \values_reg[14][6]  (.Q (\values[14] [6] ), .CK (n_121_11), .D (sps__n117));
DFF_X1 \values_reg[14][7]  (.Q (\values[14] [7] ), .CK (n_121_11), .D (spc__n127));
DFF_X1 \values_reg[14][8]  (.Q (\values[14] [8] ), .CK (n_121_11), .D (sps__n97));
DFF_X1 \values_reg[14][9]  (.Q (\values[14] [9] ), .CK (n_121_11), .D (sps__n108));
DFF_X1 \values_reg[14][10]  (.Q (\values[14] [10] ), .CK (n_121_11), .D (sps__n1));
DFF_X1 \values_reg[14][11]  (.Q (\values[14] [11] ), .CK (n_121_11), .D (sps__n11));
DFF_X1 \values_reg[14][12]  (.Q (\values[14] [12] ), .CK (n_121_11), .D (sps__n57));
DFF_X1 \values_reg[14][13]  (.Q (\values[14] [13] ), .CK (n_121_11), .D (sps__n39));
DFF_X1 \values_reg[14][14]  (.Q (\values[14] [14] ), .CK (n_121_11), .D (sps__n25));
DFF_X1 \values_reg[14][15]  (.Q (\values[14] [15] ), .CK (n_121_11), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[14]_reg  (.GCK (n_121_11), .CK (clk), .E (n_14), .SE (1'b0 ));
DFF_X1 \values_reg[13][0]  (.Q (\values[13] [0] ), .CK (n_121_10), .D (sps__n5));
DFF_X1 \values_reg[13][1]  (.Q (\values[13] [1] ), .CK (n_121_10), .D (sps__n71));
DFF_X1 \values_reg[13][2]  (.Q (\values[13] [2] ), .CK (n_121_10), .D (spc__n159));
DFF_X1 \values_reg[13][3]  (.Q (\values[13] [3] ), .CK (n_121_10), .D (sps__n77));
DFF_X1 \values_reg[13][4]  (.Q (\values[13] [4] ), .CK (n_121_10), .D (sps__n90));
DFF_X1 \values_reg[13][5]  (.Q (\values[13] [5] ), .CK (n_121_10), .D (spc__n132));
DFF_X1 \values_reg[13][6]  (.Q (\values[13] [6] ), .CK (n_121_10), .D (sps__n117));
DFF_X1 \values_reg[13][7]  (.Q (\values[13] [7] ), .CK (n_121_10), .D (spc__n127));
DFF_X1 \values_reg[13][8]  (.Q (\values[13] [8] ), .CK (n_121_10), .D (sps__n97));
DFF_X1 \values_reg[13][9]  (.Q (\values[13] [9] ), .CK (n_121_10), .D (sps__n108));
DFF_X1 \values_reg[13][10]  (.Q (\values[13] [10] ), .CK (n_121_10), .D (sps__n1));
DFF_X1 \values_reg[13][11]  (.Q (\values[13] [11] ), .CK (n_121_10), .D (sps__n12));
DFF_X1 \values_reg[13][12]  (.Q (\values[13] [12] ), .CK (n_121_10), .D (sps__n57));
DFF_X1 \values_reg[13][13]  (.Q (\values[13] [13] ), .CK (n_121_10), .D (sps__n40));
DFF_X1 \values_reg[13][14]  (.Q (\values[13] [14] ), .CK (n_121_10), .D (sps__n25));
DFF_X1 \values_reg[13][15]  (.Q (\values[13] [15] ), .CK (n_121_10), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[13]_reg  (.GCK (n_121_10), .CK (clk), .E (n_13), .SE (1'b0 ));
DFF_X1 \values_reg[12][0]  (.Q (\values[12] [0] ), .CK (n_121_9), .D (sps__n5));
DFF_X1 \values_reg[12][1]  (.Q (\values[12] [1] ), .CK (n_121_9), .D (sps__n71));
DFF_X1 \values_reg[12][2]  (.Q (\values[12] [2] ), .CK (n_121_9), .D (spc__n159));
DFF_X1 \values_reg[12][3]  (.Q (\values[12] [3] ), .CK (n_121_9), .D (sps__n77));
DFF_X1 \values_reg[12][4]  (.Q (\values[12] [4] ), .CK (n_121_9), .D (sps__n90));
DFF_X1 \values_reg[12][5]  (.Q (\values[12] [5] ), .CK (n_121_9), .D (spc__n132));
DFF_X1 \values_reg[12][6]  (.Q (\values[12] [6] ), .CK (n_121_9), .D (sps__n117));
DFF_X1 \values_reg[12][7]  (.Q (\values[12] [7] ), .CK (n_121_9), .D (spc__n127));
DFF_X1 \values_reg[12][8]  (.Q (\values[12] [8] ), .CK (n_121_9), .D (sps__n97));
DFF_X1 \values_reg[12][9]  (.Q (\values[12] [9] ), .CK (n_121_9), .D (sps__n108));
DFF_X1 \values_reg[12][10]  (.Q (\values[12] [10] ), .CK (n_121_9), .D (sps__n1));
DFF_X1 \values_reg[12][11]  (.Q (\values[12] [11] ), .CK (n_121_9), .D (sps__n11));
DFF_X1 \values_reg[12][12]  (.Q (\values[12] [12] ), .CK (n_121_9), .D (sps__n57));
DFF_X1 \values_reg[12][13]  (.Q (\values[12] [13] ), .CK (n_121_9), .D (sps__n39));
DFF_X1 \values_reg[12][14]  (.Q (\values[12] [14] ), .CK (n_121_9), .D (sps__n25));
DFF_X1 \values_reg[12][15]  (.Q (\values[12] [15] ), .CK (n_121_9), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[12]_reg  (.GCK (n_121_9), .CK (clk), .E (n_12), .SE (1'b0 ));
DFF_X1 \values_reg[11][0]  (.Q (\values[11] [0] ), .CK (n_121_8), .D (sps__n5));
DFF_X1 \values_reg[11][1]  (.Q (\values[11] [1] ), .CK (n_121_8), .D (sps__n71));
DFF_X1 \values_reg[11][2]  (.Q (\values[11] [2] ), .CK (n_121_8), .D (spc__n158));
DFF_X1 \values_reg[11][3]  (.Q (\values[11] [3] ), .CK (n_121_8), .D (sps__n77));
DFF_X1 \values_reg[11][4]  (.Q (\values[11] [4] ), .CK (n_121_8), .D (sps__n90));
DFF_X1 \values_reg[11][5]  (.Q (\values[11] [5] ), .CK (n_121_8), .D (spc__n132));
DFF_X1 \values_reg[11][6]  (.Q (\values[11] [6] ), .CK (n_121_8), .D (sps__n117));
DFF_X1 \values_reg[11][7]  (.Q (\values[11] [7] ), .CK (n_121_8), .D (spc__n127));
DFF_X1 \values_reg[11][8]  (.Q (\values[11] [8] ), .CK (n_121_8), .D (sps__n97));
DFF_X1 \values_reg[11][9]  (.Q (\values[11] [9] ), .CK (n_121_8), .D (sps__n110));
DFF_X1 \values_reg[11][10]  (.Q (\values[11] [10] ), .CK (n_121_8), .D (sps__n1));
DFF_X1 \values_reg[11][11]  (.Q (\values[11] [11] ), .CK (n_121_8), .D (sps__n11));
DFF_X1 \values_reg[11][12]  (.Q (\values[11] [12] ), .CK (n_121_8), .D (sps__n52));
DFF_X1 \values_reg[11][13]  (.Q (\values[11] [13] ), .CK (n_121_8), .D (sps__n38));
DFF_X1 \values_reg[11][14]  (.Q (\values[11] [14] ), .CK (n_121_8), .D (sps__n25));
DFF_X1 \values_reg[11][15]  (.Q (\values[11] [15] ), .CK (n_121_8), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[11]_reg  (.GCK (n_121_8), .CK (clk), .E (n_11), .SE (1'b0 ));
DFF_X1 \values_reg[10][0]  (.Q (\values[10] [0] ), .CK (n_121_7), .D (sps__n5));
DFF_X1 \values_reg[10][1]  (.Q (\values[10] [1] ), .CK (n_121_7), .D (sps__n71));
DFF_X1 \values_reg[10][2]  (.Q (\values[10] [2] ), .CK (n_121_7), .D (spc__n159));
DFF_X1 \values_reg[10][3]  (.Q (\values[10] [3] ), .CK (n_121_7), .D (sps__n77));
DFF_X1 \values_reg[10][4]  (.Q (\values[10] [4] ), .CK (n_121_7), .D (sps__n90));
DFF_X1 \values_reg[10][5]  (.Q (\values[10] [5] ), .CK (n_121_7), .D (spc__n132));
DFF_X1 \values_reg[10][6]  (.Q (\values[10] [6] ), .CK (n_121_7), .D (sps__n117));
DFF_X1 \values_reg[10][7]  (.Q (\values[10] [7] ), .CK (n_121_7), .D (spc__n127));
DFF_X1 \values_reg[10][8]  (.Q (\values[10] [8] ), .CK (n_121_7), .D (sps__n97));
DFF_X1 \values_reg[10][9]  (.Q (\values[10] [9] ), .CK (n_121_7), .D (sps__n108));
DFF_X1 \values_reg[10][10]  (.Q (\values[10] [10] ), .CK (n_121_7), .D (sps__n1));
DFF_X1 \values_reg[10][11]  (.Q (\values[10] [11] ), .CK (n_121_7), .D (sps__n11));
DFF_X1 \values_reg[10][12]  (.Q (\values[10] [12] ), .CK (n_121_7), .D (sps__n57));
DFF_X1 \values_reg[10][13]  (.Q (\values[10] [13] ), .CK (n_121_7), .D (sps__n39));
DFF_X1 \values_reg[10][14]  (.Q (\values[10] [14] ), .CK (n_121_7), .D (sps__n25));
DFF_X1 \values_reg[10][15]  (.Q (\values[10] [15] ), .CK (n_121_7), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[10]_reg  (.GCK (n_121_7), .CK (clk), .E (n_10), .SE (1'b0 ));
DFF_X1 \values_reg[9][0]  (.Q (\values[9] [0] ), .CK (n_121_6), .D (sps__n5));
DFF_X1 \values_reg[9][1]  (.Q (\values[9] [1] ), .CK (n_121_6), .D (sps__n71));
DFF_X1 \values_reg[9][2]  (.Q (\values[9] [2] ), .CK (n_121_6), .D (spc__n159));
DFF_X1 \values_reg[9][3]  (.Q (\values[9] [3] ), .CK (n_121_6), .D (sps__n77));
DFF_X1 \values_reg[9][4]  (.Q (\values[9] [4] ), .CK (n_121_6), .D (sps__n89));
DFF_X1 \values_reg[9][5]  (.Q (\values[9] [5] ), .CK (n_121_6), .D (spc__n132));
DFF_X1 \values_reg[9][6]  (.Q (\values[9] [6] ), .CK (n_121_6), .D (sps__n117));
DFF_X1 \values_reg[9][7]  (.Q (\values[9] [7] ), .CK (n_121_6), .D (spc__n127));
DFF_X1 \values_reg[9][8]  (.Q (\values[9] [8] ), .CK (n_121_6), .D (sps__n97));
DFF_X1 \values_reg[9][9]  (.Q (\values[9] [9] ), .CK (n_121_6), .D (sps__n109));
DFF_X1 \values_reg[9][10]  (.Q (\values[9] [10] ), .CK (n_121_6), .D (sps__n1));
DFF_X1 \values_reg[9][11]  (.Q (\values[9] [11] ), .CK (n_121_6), .D (sps__n12));
DFF_X1 \values_reg[9][12]  (.Q (\values[9] [12] ), .CK (n_121_6), .D (sps__n57));
DFF_X1 \values_reg[9][13]  (.Q (\values[9] [13] ), .CK (n_121_6), .D (sps__n39));
DFF_X1 \values_reg[9][14]  (.Q (\values[9] [14] ), .CK (n_121_6), .D (sps__n28));
DFF_X1 \values_reg[9][15]  (.Q (\values[9] [15] ), .CK (n_121_6), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[9]_reg  (.GCK (n_121_6), .CK (clk), .E (n_9), .SE (1'b0 ));
DFF_X1 \values_reg[8][0]  (.Q (\values[8] [0] ), .CK (n_121_5), .D (sps__n5));
DFF_X1 \values_reg[8][1]  (.Q (\values[8] [1] ), .CK (n_121_5), .D (sps__n71));
DFF_X1 \values_reg[8][2]  (.Q (\values[8] [2] ), .CK (n_121_5), .D (spc__n159));
DFF_X1 \values_reg[8][3]  (.Q (\values[8] [3] ), .CK (n_121_5), .D (sps__n77));
DFF_X1 \values_reg[8][4]  (.Q (\values[8] [4] ), .CK (n_121_5), .D (sps__n89));
DFF_X1 \values_reg[8][5]  (.Q (\values[8] [5] ), .CK (n_121_5), .D (spc__n132));
DFF_X1 \values_reg[8][6]  (.Q (\values[8] [6] ), .CK (n_121_5), .D (sps__n119));
DFF_X1 \values_reg[8][7]  (.Q (\values[8] [7] ), .CK (n_121_5), .D (spc__n127));
DFF_X1 \values_reg[8][8]  (.Q (\values[8] [8] ), .CK (n_121_5), .D (sps__n97));
DFF_X1 \values_reg[8][9]  (.Q (\values[8] [9] ), .CK (n_121_5), .D (sps__n109));
DFF_X1 \values_reg[8][10]  (.Q (\values[8] [10] ), .CK (n_121_5), .D (sps__n1));
DFF_X1 \values_reg[8][11]  (.Q (\values[8] [11] ), .CK (n_121_5), .D (sps__n12));
DFF_X1 \values_reg[8][12]  (.Q (\values[8] [12] ), .CK (n_121_5), .D (sps__n57));
DFF_X1 \values_reg[8][13]  (.Q (\values[8] [13] ), .CK (n_121_5), .D (sps__n39));
DFF_X1 \values_reg[8][14]  (.Q (\values[8] [14] ), .CK (n_121_5), .D (sps__n28));
DFF_X1 \values_reg[8][15]  (.Q (\values[8] [15] ), .CK (n_121_5), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[8]_reg  (.GCK (n_121_5), .CK (clk), .E (n_8), .SE (1'b0 ));
DFF_X1 \values_reg[7][0]  (.Q (\values[7] [0] ), .CK (n_121_4), .D (sps__n5));
DFF_X1 \values_reg[7][1]  (.Q (\values[7] [1] ), .CK (n_121_4), .D (sps__n71));
DFF_X1 \values_reg[7][2]  (.Q (\values[7] [2] ), .CK (n_121_4), .D (spc__n159));
DFF_X1 \values_reg[7][3]  (.Q (\values[7] [3] ), .CK (n_121_4), .D (sps__n77));
DFF_X1 \values_reg[7][4]  (.Q (\values[7] [4] ), .CK (n_121_4), .D (sps__n89));
DFF_X1 \values_reg[7][5]  (.Q (\values[7] [5] ), .CK (n_121_4), .D (spc__n132));
DFF_X1 \values_reg[7][6]  (.Q (\values[7] [6] ), .CK (n_121_4), .D (sps__n117));
DFF_X1 \values_reg[7][7]  (.Q (\values[7] [7] ), .CK (n_121_4), .D (spc__n127));
DFF_X1 \values_reg[7][8]  (.Q (\values[7] [8] ), .CK (n_121_4), .D (sps__n97));
DFF_X1 \values_reg[7][9]  (.Q (\values[7] [9] ), .CK (n_121_4), .D (sps__n109));
DFF_X1 \values_reg[7][10]  (.Q (\values[7] [10] ), .CK (n_121_4), .D (sps__n1));
DFF_X1 \values_reg[7][11]  (.Q (\values[7] [11] ), .CK (n_121_4), .D (sps__n12));
DFF_X1 \values_reg[7][12]  (.Q (\values[7] [12] ), .CK (n_121_4), .D (sps__n54));
DFF_X1 \values_reg[7][13]  (.Q (\values[7] [13] ), .CK (n_121_4), .D (sps__n40));
DFF_X1 \values_reg[7][14]  (.Q (\values[7] [14] ), .CK (n_121_4), .D (sps__n28));
DFF_X1 \values_reg[7][15]  (.Q (\values[7] [15] ), .CK (n_121_4), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[7]_reg  (.GCK (n_121_4), .CK (clk), .E (n_7), .SE (1'b0 ));
DFF_X1 \values_reg[6][0]  (.Q (\values[6] [0] ), .CK (n_121_3), .D (sps__n5));
DFF_X1 \values_reg[6][1]  (.Q (\values[6] [1] ), .CK (n_121_3), .D (sps__n71));
DFF_X1 \values_reg[6][2]  (.Q (\values[6] [2] ), .CK (n_121_3), .D (spc__n159));
DFF_X1 \values_reg[6][3]  (.Q (\values[6] [3] ), .CK (n_121_3), .D (sps__n77));
DFF_X1 \values_reg[6][4]  (.Q (\values[6] [4] ), .CK (n_121_3), .D (sps__n89));
DFF_X1 \values_reg[6][5]  (.Q (\values[6] [5] ), .CK (n_121_3), .D (spc__n132));
DFF_X1 \values_reg[6][6]  (.Q (\values[6] [6] ), .CK (n_121_3), .D (sps__n118));
DFF_X1 \values_reg[6][7]  (.Q (\values[6] [7] ), .CK (n_121_3), .D (spc__n127));
DFF_X1 \values_reg[6][8]  (.Q (\values[6] [8] ), .CK (n_121_3), .D (sps__n97));
DFF_X1 \values_reg[6][9]  (.Q (\values[6] [9] ), .CK (n_121_3), .D (sps__n109));
DFF_X1 \values_reg[6][10]  (.Q (\values[6] [10] ), .CK (n_121_3), .D (sps__n1));
DFF_X1 \values_reg[6][11]  (.Q (\values[6] [11] ), .CK (n_121_3), .D (sps__n12));
DFF_X1 \values_reg[6][12]  (.Q (\values[6] [12] ), .CK (n_121_3), .D (sps__n54));
DFF_X1 \values_reg[6][13]  (.Q (\values[6] [13] ), .CK (n_121_3), .D (sps__n40));
DFF_X1 \values_reg[6][14]  (.Q (\values[6] [14] ), .CK (n_121_3), .D (sps__n28));
DFF_X1 \values_reg[6][15]  (.Q (\values[6] [15] ), .CK (n_121_3), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[6]_reg  (.GCK (n_121_3), .CK (clk), .E (n_6), .SE (1'b0 ));
DFF_X1 \values_reg[5][0]  (.Q (\values[5] [0] ), .CK (n_121_2), .D (sps__n5));
DFF_X1 \values_reg[5][1]  (.Q (\values[5] [1] ), .CK (n_121_2), .D (sps__n71));
DFF_X1 \values_reg[5][2]  (.Q (\values[5] [2] ), .CK (n_121_2), .D (spc__n159));
DFF_X1 \values_reg[5][3]  (.Q (\values[5] [3] ), .CK (n_121_2), .D (sps__n77));
DFF_X1 \values_reg[5][4]  (.Q (\values[5] [4] ), .CK (n_121_2), .D (sps__n89));
DFF_X1 \values_reg[5][5]  (.Q (\values[5] [5] ), .CK (n_121_2), .D (spc__n132));
DFF_X1 \values_reg[5][6]  (.Q (\values[5] [6] ), .CK (n_121_2), .D (sps__n117));
DFF_X1 \values_reg[5][7]  (.Q (\values[5] [7] ), .CK (n_121_2), .D (spc__n127));
DFF_X1 \values_reg[5][8]  (.Q (\values[5] [8] ), .CK (n_121_2), .D (sps__n97));
DFF_X1 \values_reg[5][9]  (.Q (\values[5] [9] ), .CK (n_121_2), .D (sps__n109));
DFF_X1 \values_reg[5][10]  (.Q (\values[5] [10] ), .CK (n_121_2), .D (sps__n1));
DFF_X1 \values_reg[5][11]  (.Q (\values[5] [11] ), .CK (n_121_2), .D (sps__n12));
DFF_X1 \values_reg[5][12]  (.Q (\values[5] [12] ), .CK (n_121_2), .D (sps__n54));
DFF_X1 \values_reg[5][13]  (.Q (\values[5] [13] ), .CK (n_121_2), .D (sps__n40));
DFF_X1 \values_reg[5][14]  (.Q (\values[5] [14] ), .CK (n_121_2), .D (sps__n28));
DFF_X1 \values_reg[5][15]  (.Q (\values[5] [15] ), .CK (n_121_2), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[5]_reg  (.GCK (n_121_2), .CK (clk), .E (n_5), .SE (1'b0 ));
DFF_X1 \values_reg[4][0]  (.Q (\values[4] [0] ), .CK (n_121_1), .D (sps__n5));
DFF_X1 \values_reg[4][1]  (.Q (\values[4] [1] ), .CK (n_121_1), .D (sps__n71));
DFF_X1 \values_reg[4][2]  (.Q (\values[4] [2] ), .CK (n_121_1), .D (spc__n159));
DFF_X1 \values_reg[4][3]  (.Q (\values[4] [3] ), .CK (n_121_1), .D (sps__n77));
DFF_X1 \values_reg[4][4]  (.Q (\values[4] [4] ), .CK (n_121_1), .D (sps__n89));
DFF_X1 \values_reg[4][5]  (.Q (\values[4] [5] ), .CK (n_121_1), .D (spc__n132));
DFF_X1 \values_reg[4][6]  (.Q (\values[4] [6] ), .CK (n_121_1), .D (sps__n117));
DFF_X1 \values_reg[4][7]  (.Q (\values[4] [7] ), .CK (n_121_1), .D (spc__n127));
DFF_X1 \values_reg[4][8]  (.Q (\values[4] [8] ), .CK (n_121_1), .D (sps__n97));
DFF_X1 \values_reg[4][9]  (.Q (\values[4] [9] ), .CK (n_121_1), .D (sps__n109));
DFF_X1 \values_reg[4][10]  (.Q (\values[4] [10] ), .CK (n_121_1), .D (sps__n1));
DFF_X1 \values_reg[4][11]  (.Q (\values[4] [11] ), .CK (n_121_1), .D (sps__n12));
DFF_X1 \values_reg[4][12]  (.Q (\values[4] [12] ), .CK (n_121_1), .D (sps__n54));
DFF_X1 \values_reg[4][13]  (.Q (\values[4] [13] ), .CK (n_121_1), .D (sps__n40));
DFF_X1 \values_reg[4][14]  (.Q (\values[4] [14] ), .CK (n_121_1), .D (sps__n28));
DFF_X1 \values_reg[4][15]  (.Q (\values[4] [15] ), .CK (n_121_1), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[4]_reg  (.GCK (n_121_1), .CK (clk), .E (n_4), .SE (1'b0 ));
DFF_X1 \values_reg[3][0]  (.Q (\values[3] [0] ), .CK (n_121_0), .D (sps__n5));
DFF_X1 \values_reg[3][1]  (.Q (\values[3] [1] ), .CK (n_121_0), .D (sps__n71));
DFF_X1 \values_reg[3][2]  (.Q (\values[3] [2] ), .CK (n_121_0), .D (spc__n159));
DFF_X1 \values_reg[3][3]  (.Q (\values[3] [3] ), .CK (n_121_0), .D (sps__n77));
DFF_X1 \values_reg[3][4]  (.Q (\values[3] [4] ), .CK (n_121_0), .D (sps__n89));
DFF_X1 \values_reg[3][5]  (.Q (\values[3] [5] ), .CK (n_121_0), .D (spc__n132));
DFF_X1 \values_reg[3][6]  (.Q (\values[3] [6] ), .CK (n_121_0), .D (sps__n118));
DFF_X1 \values_reg[3][7]  (.Q (\values[3] [7] ), .CK (n_121_0), .D (spc__n127));
DFF_X1 \values_reg[3][8]  (.Q (\values[3] [8] ), .CK (n_121_0), .D (sps__n97));
DFF_X1 \values_reg[3][9]  (.Q (\values[3] [9] ), .CK (n_121_0), .D (sps__n109));
DFF_X1 \values_reg[3][10]  (.Q (\values[3] [10] ), .CK (n_121_0), .D (sps__n1));
DFF_X1 \values_reg[3][11]  (.Q (\values[3] [11] ), .CK (n_121_0), .D (sps__n12));
DFF_X1 \values_reg[3][12]  (.Q (\values[3] [12] ), .CK (n_121_0), .D (sps__n54));
DFF_X1 \values_reg[3][13]  (.Q (\values[3] [13] ), .CK (n_121_0), .D (sps__n40));
DFF_X1 \values_reg[3][14]  (.Q (\values[3] [14] ), .CK (n_121_0), .D (sps__n28));
DFF_X1 \values_reg[3][15]  (.Q (\values[3] [15] ), .CK (n_121_0), .D (sps__n49));
CLKGATETST_X1 \clk_gate_values_reg[3]_reg  (.GCK (n_121_0), .CK (clk), .E (n_3), .SE (1'b0 ));
BUF_X16 sps__L1_c1 (.Z (sps__n1), .A (\values[10] ));
INV_X4 sps__L1_c4 (.ZN (sps__n4), .A (\values[0] ));
INV_X16 sps__L2_c5 (.ZN (sps__n5), .A (sps__n4));
BUF_X4 sps__L1_c10 (.Z (sps__n10), .A (\values[11] ));
CLKBUF_X3 sps__L2_c11 (.Z (sps__n11), .A (sps__n10));
BUF_X8 sps__L2_c12 (.Z (sps__n12), .A (sps__n10));
BUF_X8 spc__L1_c157 (.Z (spc__n157), .A (\values[2] ));
CLKBUF_X3 sps__L2_c14 (.Z (sps__n14), .A (sps__n10));
BUF_X4 sps__L1_c25 (.Z (sps__n25), .A (\values[14] ));
CLKBUF_X3 spc__L1_c158 (.Z (spc__n158), .A (\values[2] ));
BUF_X2 sps__L2_c27 (.Z (sps__n27), .A (sps__n25));
BUF_X16 sps__L2_c28 (.Z (sps__n28), .A (sps__n25));
BUF_X4 sps__L1_c37 (.Z (sps__n37), .A (\values[13] ));
CLKBUF_X3 sps__L2_c38 (.Z (sps__n38), .A (sps__n37));
BUF_X1 sps__L2_c39 (.Z (sps__n39), .A (sps__n37));
BUF_X16 sps__L2_c40 (.Z (sps__n40), .A (sps__n37));
BUF_X16 sps__L1_c49 (.Z (sps__n49), .A (\values[15] ));
BUF_X4 sps__L1_c52 (.Z (sps__n52), .A (\values[12] ));
BUF_X8 spc__L1_c159 (.Z (spc__n159), .A (\values[2] ));
BUF_X4 sps__L2_c54 (.Z (sps__n54), .A (sps__n52));
BUF_X8 sps__L2_c55 (.Z (sps__n55), .A (sps__n52));
BUF_X1 sps__L2_c57 (.Z (sps__n57), .A (sps__n52));
INV_X4 sps__L1_c70 (.ZN (sps__n70), .A (\values[1] ));
INV_X16 sps__L2_c71 (.ZN (sps__n71), .A (sps__n70));
BUF_X4 sps__L1_c76 (.Z (sps__n76), .A (\values[3] ));
BUF_X8 sps__L2_c77 (.Z (sps__n77), .A (sps__n76));
CLKBUF_X3 sps__L2_c78 (.Z (sps__n78), .A (sps__n76));
BUF_X8 sps__L2_c79 (.Z (sps__n79), .A (sps__n76));
BUF_X4 sps__L1_c88 (.Z (sps__n88), .A (\values[4] ));
BUF_X16 sps__L2_c89 (.Z (sps__n89), .A (sps__n88));
CLKBUF_X3 sps__L2_c90 (.Z (sps__n90), .A (sps__n88));
BUF_X16 sps__L1_c97 (.Z (sps__n97), .A (\values[8] ));
CLKBUF_X3 sps__L1_c108 (.Z (sps__n108), .A (\values[9] ));
BUF_X8 sps__L1_c109 (.Z (sps__n109), .A (\values[9] ));
CLKBUF_X3 sps__L1_c110 (.Z (sps__n110), .A (\values[9] ));
BUF_X4 sps__L1_c117 (.Z (sps__n117), .A (\values[6] ));
BUF_X8 sps__L1_c118 (.Z (sps__n118), .A (\values[6] ));
CLKBUF_X3 sps__L1_c119 (.Z (sps__n119), .A (\values[6] ));
BUF_X8 spc__L1_c126 (.Z (spc__n126), .A (\values[7] ));
BUF_X8 spc__L1_c127 (.Z (spc__n127), .A (\values[7] ));
BUF_X16 spc__L1_c132 (.Z (spc__n132), .A (\values[5] ));

endmodule //Neuron_Layer


