/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 05:33:27 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2542322260 */

module Neuron_Layer(clk, load_en, load_value, load_address, reset, \values[0] , 
      \values[1] , \values[2] , \values[3] , \values[4] , \values[5] , 
      \values[6] , \values[7] , \values[8] , \values[9] , \values[10] , 
      \values[11] , \values[12] , \values[13] , \values[14] , \values[15] , 
      \values[16] , \values[17] , \values[18] , \values[19] , \values[20] , 
      \values[21] , \values[22] , \values[23] , \values[24] , \values[25] , 
      \values[26] , \values[27] , \values[28] , \values[29] , \values[30] , 
      \values[31] , \values[32] , \values[33] , \values[34] , \values[35] , 
      \values[36] , \values[37] , \values[38] , \values[39] , \values[40] , 
      \values[41] , \values[42] , \values[43] , \values[44] , \values[45] , 
      \values[46] , \values[47] , \values[48] , \values[49] , \values[50] , 
      \values[51] , \values[52] , \values[53] , \values[54] , \values[55] , 
      \values[56] , \values[57] , \values[58] , \values[59] , \values[60] , 
      \values[61] , \values[62] , \values[63] , \values[64] , \values[65] , 
      \values[66] , \values[67] , \values[68] , \values[69] , \values[70] , 
      \values[71] , \values[72] , \values[73] , \values[74] , \values[75] , 
      \values[76] , \values[77] , \values[78] , \values[79] , \values[80] , 
      \values[81] , \values[82] , \values[83] , \values[84] , \values[85] , 
      \values[86] , \values[87] , \values[88] , \values[89] , \values[90] , 
      \values[91] , \values[92] , \values[93] , \values[94] , \values[95] , 
      \values[96] , \values[97] , \values[98] , \values[99] , \values[100] , 
      \values[101] , \values[102] , \values[103] , \values[104] , \values[105] , 
      \values[106] , \values[107] , \values[108] , \values[109] , \values[110] , 
      \values[111] , \values[112] , \values[113] , \values[114] , \values[115] , 
      \values[116] , \values[117] , \values[118] , \values[119] );
   input clk;
   input load_en;
   input [15:0]load_value;
   input [15:0]load_address;
   input reset;
   output [15:0]\values[0] ;
   output [15:0]\values[1] ;
   output [15:0]\values[2] ;
   output [15:0]\values[3] ;
   output [15:0]\values[4] ;
   output [15:0]\values[5] ;
   output [15:0]\values[6] ;
   output [15:0]\values[7] ;
   output [15:0]\values[8] ;
   output [15:0]\values[9] ;
   output [15:0]\values[10] ;
   output [15:0]\values[11] ;
   output [15:0]\values[12] ;
   output [15:0]\values[13] ;
   output [15:0]\values[14] ;
   output [15:0]\values[15] ;
   output [15:0]\values[16] ;
   output [15:0]\values[17] ;
   output [15:0]\values[18] ;
   output [15:0]\values[19] ;
   output [15:0]\values[20] ;
   output [15:0]\values[21] ;
   output [15:0]\values[22] ;
   output [15:0]\values[23] ;
   output [15:0]\values[24] ;
   output [15:0]\values[25] ;
   output [15:0]\values[26] ;
   output [15:0]\values[27] ;
   output [15:0]\values[28] ;
   output [15:0]\values[29] ;
   output [15:0]\values[30] ;
   output [15:0]\values[31] ;
   output [15:0]\values[32] ;
   output [15:0]\values[33] ;
   output [15:0]\values[34] ;
   output [15:0]\values[35] ;
   output [15:0]\values[36] ;
   output [15:0]\values[37] ;
   output [15:0]\values[38] ;
   output [15:0]\values[39] ;
   output [15:0]\values[40] ;
   output [15:0]\values[41] ;
   output [15:0]\values[42] ;
   output [15:0]\values[43] ;
   output [15:0]\values[44] ;
   output [15:0]\values[45] ;
   output [15:0]\values[46] ;
   output [15:0]\values[47] ;
   output [15:0]\values[48] ;
   output [15:0]\values[49] ;
   output [15:0]\values[50] ;
   output [15:0]\values[51] ;
   output [15:0]\values[52] ;
   output [15:0]\values[53] ;
   output [15:0]\values[54] ;
   output [15:0]\values[55] ;
   output [15:0]\values[56] ;
   output [15:0]\values[57] ;
   output [15:0]\values[58] ;
   output [15:0]\values[59] ;
   output [15:0]\values[60] ;
   output [15:0]\values[61] ;
   output [15:0]\values[62] ;
   output [15:0]\values[63] ;
   output [15:0]\values[64] ;
   output [15:0]\values[65] ;
   output [15:0]\values[66] ;
   output [15:0]\values[67] ;
   output [15:0]\values[68] ;
   output [15:0]\values[69] ;
   output [15:0]\values[70] ;
   output [15:0]\values[71] ;
   output [15:0]\values[72] ;
   output [15:0]\values[73] ;
   output [15:0]\values[74] ;
   output [15:0]\values[75] ;
   output [15:0]\values[76] ;
   output [15:0]\values[77] ;
   output [15:0]\values[78] ;
   output [15:0]\values[79] ;
   output [15:0]\values[80] ;
   output [15:0]\values[81] ;
   output [15:0]\values[82] ;
   output [15:0]\values[83] ;
   output [15:0]\values[84] ;
   output [15:0]\values[85] ;
   output [15:0]\values[86] ;
   output [15:0]\values[87] ;
   output [15:0]\values[88] ;
   output [15:0]\values[89] ;
   output [15:0]\values[90] ;
   output [15:0]\values[91] ;
   output [15:0]\values[92] ;
   output [15:0]\values[93] ;
   output [15:0]\values[94] ;
   output [15:0]\values[95] ;
   output [15:0]\values[96] ;
   output [15:0]\values[97] ;
   output [15:0]\values[98] ;
   output [15:0]\values[99] ;
   output [15:0]\values[100] ;
   output [15:0]\values[101] ;
   output [15:0]\values[102] ;
   output [15:0]\values[103] ;
   output [15:0]\values[104] ;
   output [15:0]\values[105] ;
   output [15:0]\values[106] ;
   output [15:0]\values[107] ;
   output [15:0]\values[108] ;
   output [15:0]\values[109] ;
   output [15:0]\values[110] ;
   output [15:0]\values[111] ;
   output [15:0]\values[112] ;
   output [15:0]\values[113] ;
   output [15:0]\values[114] ;
   output [15:0]\values[115] ;
   output [15:0]\values[116] ;
   output [15:0]\values[117] ;
   output [15:0]\values[118] ;
   output [15:0]\values[119] ;

   wire n_121_0;
   wire n_121_1;
   wire n_121_2;
   wire n_121_3;
   wire n_121_4;
   wire n_121_5;
   wire n_121_6;
   wire n_121_7;
   wire n_121_8;
   wire n_121_9;
   wire n_121_10;
   wire n_121_11;
   wire n_121_12;
   wire n_121_13;
   wire n_121_14;
   wire n_121_15;
   wire n_121_16;
   wire n_121_17;
   wire n_121_18;
   wire n_121_19;
   wire n_121_20;
   wire n_121_21;
   wire n_121_22;
   wire n_121_23;
   wire n_121_24;
   wire n_121_25;
   wire n_121_26;
   wire n_121_27;
   wire n_121_28;
   wire n_121_29;
   wire n_121_30;
   wire n_121_31;
   wire n_121_32;
   wire n_121_33;
   wire n_121_34;
   wire n_121_35;
   wire n_121_36;
   wire n_121_37;
   wire n_121_38;
   wire n_121_39;
   wire n_121_40;
   wire n_121_41;
   wire n_121_42;
   wire n_121_43;
   wire n_121_44;
   wire n_121_45;
   wire n_121_46;
   wire n_121_47;
   wire n_121_48;
   wire n_121_49;
   wire n_121_50;
   wire n_121_51;
   wire n_121_52;
   wire n_121_53;
   wire n_121_54;
   wire n_121_55;
   wire n_121_56;
   wire n_121_57;
   wire n_121_58;
   wire n_121_59;
   wire n_121_60;
   wire n_121_61;
   wire n_121_62;
   wire n_121_63;
   wire n_121_64;
   wire n_121_65;
   wire n_121_66;
   wire n_121_67;
   wire n_121_68;
   wire n_121_69;
   wire n_121_70;
   wire n_121_71;
   wire n_121_72;
   wire n_121_73;
   wire n_121_74;
   wire n_121_75;
   wire n_121_76;
   wire n_121_77;
   wire n_121_78;
   wire n_121_79;
   wire n_121_80;
   wire n_121_81;
   wire n_121_82;
   wire n_121_83;
   wire n_121_84;
   wire n_121_85;
   wire n_121_86;
   wire n_121_87;
   wire n_121_88;
   wire n_121_89;
   wire n_121_90;
   wire n_121_91;
   wire n_121_92;
   wire n_121_93;
   wire n_122_0;
   wire n_122_1;
   wire n_122_2;
   wire n_122_3;
   wire n_122_4;
   wire n_122_5;
   wire n_122_6;
   wire n_122_7;
   wire n_122_8;
   wire n_122_9;
   wire n_122_10;
   wire n_122_11;
   wire n_122_12;
   wire n_122_13;
   wire n_122_14;
   wire n_122_15;
   wire n_122_16;
   wire n_122_17;
   wire n_122_18;
   wire n_122_19;
   wire n_122_20;
   wire n_122_21;
   wire n_122_22;
   wire n_122_23;
   wire n_122_24;
   wire n_122_25;
   wire n_0_0_0;
   wire [15:0]values;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;

   CLKGATETST_X1 \clk_gate_values_reg[3]_reg  (.CK(clk), .E(n_3), .SE(1'b0), 
      .GCK(n_121_0));
   DFF_X1 \values_reg[3][15]  (.D(values[15]), .CK(n_121_0), .Q(\values[3] [15]), 
      .QN());
   DFF_X1 \values_reg[3][14]  (.D(values[14]), .CK(n_121_0), .Q(\values[3] [14]), 
      .QN());
   DFF_X1 \values_reg[3][13]  (.D(values[13]), .CK(n_121_0), .Q(\values[3] [13]), 
      .QN());
   DFF_X1 \values_reg[3][12]  (.D(values[12]), .CK(n_121_0), .Q(\values[3] [12]), 
      .QN());
   DFF_X1 \values_reg[3][11]  (.D(values[11]), .CK(n_121_0), .Q(\values[3] [11]), 
      .QN());
   DFF_X1 \values_reg[3][10]  (.D(values[10]), .CK(n_121_0), .Q(\values[3] [10]), 
      .QN());
   DFF_X1 \values_reg[3][9]  (.D(values[9]), .CK(n_121_0), .Q(\values[3] [9]), 
      .QN());
   DFF_X1 \values_reg[3][8]  (.D(values[8]), .CK(n_121_0), .Q(\values[3] [8]), 
      .QN());
   DFF_X1 \values_reg[3][7]  (.D(values[7]), .CK(n_121_0), .Q(\values[3] [7]), 
      .QN());
   DFF_X1 \values_reg[3][6]  (.D(values[6]), .CK(n_121_0), .Q(\values[3] [6]), 
      .QN());
   DFF_X1 \values_reg[3][5]  (.D(values[5]), .CK(n_121_0), .Q(\values[3] [5]), 
      .QN());
   DFF_X1 \values_reg[3][4]  (.D(values[4]), .CK(n_121_0), .Q(\values[3] [4]), 
      .QN());
   DFF_X1 \values_reg[3][3]  (.D(values[3]), .CK(n_121_0), .Q(\values[3] [3]), 
      .QN());
   DFF_X1 \values_reg[3][2]  (.D(values[2]), .CK(n_121_0), .Q(\values[3] [2]), 
      .QN());
   DFF_X1 \values_reg[3][1]  (.D(values[1]), .CK(n_121_0), .Q(\values[3] [1]), 
      .QN());
   DFF_X1 \values_reg[3][0]  (.D(values[0]), .CK(n_121_0), .Q(\values[3] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[4]_reg  (.CK(clk), .E(n_4), .SE(1'b0), 
      .GCK(n_121_1));
   DFF_X1 \values_reg[4][15]  (.D(values[15]), .CK(n_121_1), .Q(\values[4] [15]), 
      .QN());
   DFF_X1 \values_reg[4][14]  (.D(values[14]), .CK(n_121_1), .Q(\values[4] [14]), 
      .QN());
   DFF_X1 \values_reg[4][13]  (.D(values[13]), .CK(n_121_1), .Q(\values[4] [13]), 
      .QN());
   DFF_X1 \values_reg[4][12]  (.D(values[12]), .CK(n_121_1), .Q(\values[4] [12]), 
      .QN());
   DFF_X1 \values_reg[4][11]  (.D(values[11]), .CK(n_121_1), .Q(\values[4] [11]), 
      .QN());
   DFF_X1 \values_reg[4][10]  (.D(values[10]), .CK(n_121_1), .Q(\values[4] [10]), 
      .QN());
   DFF_X1 \values_reg[4][9]  (.D(values[9]), .CK(n_121_1), .Q(\values[4] [9]), 
      .QN());
   DFF_X1 \values_reg[4][8]  (.D(values[8]), .CK(n_121_1), .Q(\values[4] [8]), 
      .QN());
   DFF_X1 \values_reg[4][7]  (.D(values[7]), .CK(n_121_1), .Q(\values[4] [7]), 
      .QN());
   DFF_X1 \values_reg[4][6]  (.D(values[6]), .CK(n_121_1), .Q(\values[4] [6]), 
      .QN());
   DFF_X1 \values_reg[4][5]  (.D(values[5]), .CK(n_121_1), .Q(\values[4] [5]), 
      .QN());
   DFF_X1 \values_reg[4][4]  (.D(values[4]), .CK(n_121_1), .Q(\values[4] [4]), 
      .QN());
   DFF_X1 \values_reg[4][3]  (.D(values[3]), .CK(n_121_1), .Q(\values[4] [3]), 
      .QN());
   DFF_X1 \values_reg[4][2]  (.D(values[2]), .CK(n_121_1), .Q(\values[4] [2]), 
      .QN());
   DFF_X1 \values_reg[4][1]  (.D(values[1]), .CK(n_121_1), .Q(\values[4] [1]), 
      .QN());
   DFF_X1 \values_reg[4][0]  (.D(values[0]), .CK(n_121_1), .Q(\values[4] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[5]_reg  (.CK(clk), .E(n_5), .SE(1'b0), 
      .GCK(n_121_2));
   DFF_X1 \values_reg[5][15]  (.D(values[15]), .CK(n_121_2), .Q(\values[5] [15]), 
      .QN());
   DFF_X1 \values_reg[5][14]  (.D(values[14]), .CK(n_121_2), .Q(\values[5] [14]), 
      .QN());
   DFF_X1 \values_reg[5][13]  (.D(values[13]), .CK(n_121_2), .Q(\values[5] [13]), 
      .QN());
   DFF_X1 \values_reg[5][12]  (.D(values[12]), .CK(n_121_2), .Q(\values[5] [12]), 
      .QN());
   DFF_X1 \values_reg[5][11]  (.D(values[11]), .CK(n_121_2), .Q(\values[5] [11]), 
      .QN());
   DFF_X1 \values_reg[5][10]  (.D(values[10]), .CK(n_121_2), .Q(\values[5] [10]), 
      .QN());
   DFF_X1 \values_reg[5][9]  (.D(values[9]), .CK(n_121_2), .Q(\values[5] [9]), 
      .QN());
   DFF_X1 \values_reg[5][8]  (.D(values[8]), .CK(n_121_2), .Q(\values[5] [8]), 
      .QN());
   DFF_X1 \values_reg[5][7]  (.D(values[7]), .CK(n_121_2), .Q(\values[5] [7]), 
      .QN());
   DFF_X1 \values_reg[5][6]  (.D(values[6]), .CK(n_121_2), .Q(\values[5] [6]), 
      .QN());
   DFF_X1 \values_reg[5][5]  (.D(values[5]), .CK(n_121_2), .Q(\values[5] [5]), 
      .QN());
   DFF_X1 \values_reg[5][4]  (.D(values[4]), .CK(n_121_2), .Q(\values[5] [4]), 
      .QN());
   DFF_X1 \values_reg[5][3]  (.D(values[3]), .CK(n_121_2), .Q(\values[5] [3]), 
      .QN());
   DFF_X1 \values_reg[5][2]  (.D(values[2]), .CK(n_121_2), .Q(\values[5] [2]), 
      .QN());
   DFF_X1 \values_reg[5][1]  (.D(values[1]), .CK(n_121_2), .Q(\values[5] [1]), 
      .QN());
   DFF_X1 \values_reg[5][0]  (.D(values[0]), .CK(n_121_2), .Q(\values[5] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[6]_reg  (.CK(clk), .E(n_6), .SE(1'b0), 
      .GCK(n_121_3));
   DFF_X1 \values_reg[6][15]  (.D(values[15]), .CK(n_121_3), .Q(\values[6] [15]), 
      .QN());
   DFF_X1 \values_reg[6][14]  (.D(values[14]), .CK(n_121_3), .Q(\values[6] [14]), 
      .QN());
   DFF_X1 \values_reg[6][13]  (.D(values[13]), .CK(n_121_3), .Q(\values[6] [13]), 
      .QN());
   DFF_X1 \values_reg[6][12]  (.D(values[12]), .CK(n_121_3), .Q(\values[6] [12]), 
      .QN());
   DFF_X1 \values_reg[6][11]  (.D(values[11]), .CK(n_121_3), .Q(\values[6] [11]), 
      .QN());
   DFF_X1 \values_reg[6][10]  (.D(values[10]), .CK(n_121_3), .Q(\values[6] [10]), 
      .QN());
   DFF_X1 \values_reg[6][9]  (.D(values[9]), .CK(n_121_3), .Q(\values[6] [9]), 
      .QN());
   DFF_X1 \values_reg[6][8]  (.D(values[8]), .CK(n_121_3), .Q(\values[6] [8]), 
      .QN());
   DFF_X1 \values_reg[6][7]  (.D(values[7]), .CK(n_121_3), .Q(\values[6] [7]), 
      .QN());
   DFF_X1 \values_reg[6][6]  (.D(values[6]), .CK(n_121_3), .Q(\values[6] [6]), 
      .QN());
   DFF_X1 \values_reg[6][5]  (.D(values[5]), .CK(n_121_3), .Q(\values[6] [5]), 
      .QN());
   DFF_X1 \values_reg[6][4]  (.D(values[4]), .CK(n_121_3), .Q(\values[6] [4]), 
      .QN());
   DFF_X1 \values_reg[6][3]  (.D(values[3]), .CK(n_121_3), .Q(\values[6] [3]), 
      .QN());
   DFF_X1 \values_reg[6][2]  (.D(values[2]), .CK(n_121_3), .Q(\values[6] [2]), 
      .QN());
   DFF_X1 \values_reg[6][1]  (.D(values[1]), .CK(n_121_3), .Q(\values[6] [1]), 
      .QN());
   DFF_X1 \values_reg[6][0]  (.D(values[0]), .CK(n_121_3), .Q(\values[6] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[7]_reg  (.CK(clk), .E(n_7), .SE(1'b0), 
      .GCK(n_121_4));
   DFF_X1 \values_reg[7][15]  (.D(values[15]), .CK(n_121_4), .Q(\values[7] [15]), 
      .QN());
   DFF_X1 \values_reg[7][14]  (.D(values[14]), .CK(n_121_4), .Q(\values[7] [14]), 
      .QN());
   DFF_X1 \values_reg[7][13]  (.D(values[13]), .CK(n_121_4), .Q(\values[7] [13]), 
      .QN());
   DFF_X1 \values_reg[7][12]  (.D(values[12]), .CK(n_121_4), .Q(\values[7] [12]), 
      .QN());
   DFF_X1 \values_reg[7][11]  (.D(values[11]), .CK(n_121_4), .Q(\values[7] [11]), 
      .QN());
   DFF_X1 \values_reg[7][10]  (.D(values[10]), .CK(n_121_4), .Q(\values[7] [10]), 
      .QN());
   DFF_X1 \values_reg[7][9]  (.D(values[9]), .CK(n_121_4), .Q(\values[7] [9]), 
      .QN());
   DFF_X1 \values_reg[7][8]  (.D(values[8]), .CK(n_121_4), .Q(\values[7] [8]), 
      .QN());
   DFF_X1 \values_reg[7][7]  (.D(values[7]), .CK(n_121_4), .Q(\values[7] [7]), 
      .QN());
   DFF_X1 \values_reg[7][6]  (.D(values[6]), .CK(n_121_4), .Q(\values[7] [6]), 
      .QN());
   DFF_X1 \values_reg[7][5]  (.D(values[5]), .CK(n_121_4), .Q(\values[7] [5]), 
      .QN());
   DFF_X1 \values_reg[7][4]  (.D(values[4]), .CK(n_121_4), .Q(\values[7] [4]), 
      .QN());
   DFF_X1 \values_reg[7][3]  (.D(values[3]), .CK(n_121_4), .Q(\values[7] [3]), 
      .QN());
   DFF_X1 \values_reg[7][2]  (.D(values[2]), .CK(n_121_4), .Q(\values[7] [2]), 
      .QN());
   DFF_X1 \values_reg[7][1]  (.D(values[1]), .CK(n_121_4), .Q(\values[7] [1]), 
      .QN());
   DFF_X1 \values_reg[7][0]  (.D(values[0]), .CK(n_121_4), .Q(\values[7] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[8]_reg  (.CK(clk), .E(n_8), .SE(1'b0), 
      .GCK(n_121_5));
   DFF_X1 \values_reg[8][15]  (.D(values[15]), .CK(n_121_5), .Q(\values[8] [15]), 
      .QN());
   DFF_X1 \values_reg[8][14]  (.D(values[14]), .CK(n_121_5), .Q(\values[8] [14]), 
      .QN());
   DFF_X1 \values_reg[8][13]  (.D(values[13]), .CK(n_121_5), .Q(\values[8] [13]), 
      .QN());
   DFF_X1 \values_reg[8][12]  (.D(values[12]), .CK(n_121_5), .Q(\values[8] [12]), 
      .QN());
   DFF_X1 \values_reg[8][11]  (.D(values[11]), .CK(n_121_5), .Q(\values[8] [11]), 
      .QN());
   DFF_X1 \values_reg[8][10]  (.D(values[10]), .CK(n_121_5), .Q(\values[8] [10]), 
      .QN());
   DFF_X1 \values_reg[8][9]  (.D(values[9]), .CK(n_121_5), .Q(\values[8] [9]), 
      .QN());
   DFF_X1 \values_reg[8][8]  (.D(values[8]), .CK(n_121_5), .Q(\values[8] [8]), 
      .QN());
   DFF_X1 \values_reg[8][7]  (.D(values[7]), .CK(n_121_5), .Q(\values[8] [7]), 
      .QN());
   DFF_X1 \values_reg[8][6]  (.D(values[6]), .CK(n_121_5), .Q(\values[8] [6]), 
      .QN());
   DFF_X1 \values_reg[8][5]  (.D(values[5]), .CK(n_121_5), .Q(\values[8] [5]), 
      .QN());
   DFF_X1 \values_reg[8][4]  (.D(values[4]), .CK(n_121_5), .Q(\values[8] [4]), 
      .QN());
   DFF_X1 \values_reg[8][3]  (.D(values[3]), .CK(n_121_5), .Q(\values[8] [3]), 
      .QN());
   DFF_X1 \values_reg[8][2]  (.D(values[2]), .CK(n_121_5), .Q(\values[8] [2]), 
      .QN());
   DFF_X1 \values_reg[8][1]  (.D(values[1]), .CK(n_121_5), .Q(\values[8] [1]), 
      .QN());
   DFF_X1 \values_reg[8][0]  (.D(values[0]), .CK(n_121_5), .Q(\values[8] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[9]_reg  (.CK(clk), .E(n_9), .SE(1'b0), 
      .GCK(n_121_6));
   DFF_X1 \values_reg[9][15]  (.D(values[15]), .CK(n_121_6), .Q(\values[9] [15]), 
      .QN());
   DFF_X1 \values_reg[9][14]  (.D(values[14]), .CK(n_121_6), .Q(\values[9] [14]), 
      .QN());
   DFF_X1 \values_reg[9][13]  (.D(values[13]), .CK(n_121_6), .Q(\values[9] [13]), 
      .QN());
   DFF_X1 \values_reg[9][12]  (.D(values[12]), .CK(n_121_6), .Q(\values[9] [12]), 
      .QN());
   DFF_X1 \values_reg[9][11]  (.D(values[11]), .CK(n_121_6), .Q(\values[9] [11]), 
      .QN());
   DFF_X1 \values_reg[9][10]  (.D(values[10]), .CK(n_121_6), .Q(\values[9] [10]), 
      .QN());
   DFF_X1 \values_reg[9][9]  (.D(values[9]), .CK(n_121_6), .Q(\values[9] [9]), 
      .QN());
   DFF_X1 \values_reg[9][8]  (.D(values[8]), .CK(n_121_6), .Q(\values[9] [8]), 
      .QN());
   DFF_X1 \values_reg[9][7]  (.D(values[7]), .CK(n_121_6), .Q(\values[9] [7]), 
      .QN());
   DFF_X1 \values_reg[9][6]  (.D(values[6]), .CK(n_121_6), .Q(\values[9] [6]), 
      .QN());
   DFF_X1 \values_reg[9][5]  (.D(values[5]), .CK(n_121_6), .Q(\values[9] [5]), 
      .QN());
   DFF_X1 \values_reg[9][4]  (.D(values[4]), .CK(n_121_6), .Q(\values[9] [4]), 
      .QN());
   DFF_X1 \values_reg[9][3]  (.D(values[3]), .CK(n_121_6), .Q(\values[9] [3]), 
      .QN());
   DFF_X1 \values_reg[9][2]  (.D(values[2]), .CK(n_121_6), .Q(\values[9] [2]), 
      .QN());
   DFF_X1 \values_reg[9][1]  (.D(values[1]), .CK(n_121_6), .Q(\values[9] [1]), 
      .QN());
   DFF_X1 \values_reg[9][0]  (.D(values[0]), .CK(n_121_6), .Q(\values[9] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[10]_reg  (.CK(clk), .E(n_10), .SE(1'b0), 
      .GCK(n_121_7));
   DFF_X1 \values_reg[10][15]  (.D(values[15]), .CK(n_121_7), .Q(
      \values[10] [15]), .QN());
   DFF_X1 \values_reg[10][14]  (.D(values[14]), .CK(n_121_7), .Q(
      \values[10] [14]), .QN());
   DFF_X1 \values_reg[10][13]  (.D(values[13]), .CK(n_121_7), .Q(
      \values[10] [13]), .QN());
   DFF_X1 \values_reg[10][12]  (.D(values[12]), .CK(n_121_7), .Q(
      \values[10] [12]), .QN());
   DFF_X1 \values_reg[10][11]  (.D(values[11]), .CK(n_121_7), .Q(
      \values[10] [11]), .QN());
   DFF_X1 \values_reg[10][10]  (.D(values[10]), .CK(n_121_7), .Q(
      \values[10] [10]), .QN());
   DFF_X1 \values_reg[10][9]  (.D(values[9]), .CK(n_121_7), .Q(\values[10] [9]), 
      .QN());
   DFF_X1 \values_reg[10][8]  (.D(values[8]), .CK(n_121_7), .Q(\values[10] [8]), 
      .QN());
   DFF_X1 \values_reg[10][7]  (.D(values[7]), .CK(n_121_7), .Q(\values[10] [7]), 
      .QN());
   DFF_X1 \values_reg[10][6]  (.D(values[6]), .CK(n_121_7), .Q(\values[10] [6]), 
      .QN());
   DFF_X1 \values_reg[10][5]  (.D(values[5]), .CK(n_121_7), .Q(\values[10] [5]), 
      .QN());
   DFF_X1 \values_reg[10][4]  (.D(values[4]), .CK(n_121_7), .Q(\values[10] [4]), 
      .QN());
   DFF_X1 \values_reg[10][3]  (.D(values[3]), .CK(n_121_7), .Q(\values[10] [3]), 
      .QN());
   DFF_X1 \values_reg[10][2]  (.D(values[2]), .CK(n_121_7), .Q(\values[10] [2]), 
      .QN());
   DFF_X1 \values_reg[10][1]  (.D(values[1]), .CK(n_121_7), .Q(\values[10] [1]), 
      .QN());
   DFF_X1 \values_reg[10][0]  (.D(values[0]), .CK(n_121_7), .Q(\values[10] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[11]_reg  (.CK(clk), .E(n_11), .SE(1'b0), 
      .GCK(n_121_8));
   DFF_X1 \values_reg[11][15]  (.D(values[15]), .CK(n_121_8), .Q(
      \values[11] [15]), .QN());
   DFF_X1 \values_reg[11][14]  (.D(values[14]), .CK(n_121_8), .Q(
      \values[11] [14]), .QN());
   DFF_X1 \values_reg[11][13]  (.D(values[13]), .CK(n_121_8), .Q(
      \values[11] [13]), .QN());
   DFF_X1 \values_reg[11][12]  (.D(values[12]), .CK(n_121_8), .Q(
      \values[11] [12]), .QN());
   DFF_X1 \values_reg[11][11]  (.D(values[11]), .CK(n_121_8), .Q(
      \values[11] [11]), .QN());
   DFF_X1 \values_reg[11][10]  (.D(values[10]), .CK(n_121_8), .Q(
      \values[11] [10]), .QN());
   DFF_X1 \values_reg[11][9]  (.D(values[9]), .CK(n_121_8), .Q(\values[11] [9]), 
      .QN());
   DFF_X1 \values_reg[11][8]  (.D(values[8]), .CK(n_121_8), .Q(\values[11] [8]), 
      .QN());
   DFF_X1 \values_reg[11][7]  (.D(values[7]), .CK(n_121_8), .Q(\values[11] [7]), 
      .QN());
   DFF_X1 \values_reg[11][6]  (.D(values[6]), .CK(n_121_8), .Q(\values[11] [6]), 
      .QN());
   DFF_X1 \values_reg[11][5]  (.D(values[5]), .CK(n_121_8), .Q(\values[11] [5]), 
      .QN());
   DFF_X1 \values_reg[11][4]  (.D(values[4]), .CK(n_121_8), .Q(\values[11] [4]), 
      .QN());
   DFF_X1 \values_reg[11][3]  (.D(values[3]), .CK(n_121_8), .Q(\values[11] [3]), 
      .QN());
   DFF_X1 \values_reg[11][2]  (.D(values[2]), .CK(n_121_8), .Q(\values[11] [2]), 
      .QN());
   DFF_X1 \values_reg[11][1]  (.D(values[1]), .CK(n_121_8), .Q(\values[11] [1]), 
      .QN());
   DFF_X1 \values_reg[11][0]  (.D(values[0]), .CK(n_121_8), .Q(\values[11] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[12]_reg  (.CK(clk), .E(n_12), .SE(1'b0), 
      .GCK(n_121_9));
   DFF_X1 \values_reg[12][15]  (.D(values[15]), .CK(n_121_9), .Q(
      \values[12] [15]), .QN());
   DFF_X1 \values_reg[12][14]  (.D(values[14]), .CK(n_121_9), .Q(
      \values[12] [14]), .QN());
   DFF_X1 \values_reg[12][13]  (.D(values[13]), .CK(n_121_9), .Q(
      \values[12] [13]), .QN());
   DFF_X1 \values_reg[12][12]  (.D(values[12]), .CK(n_121_9), .Q(
      \values[12] [12]), .QN());
   DFF_X1 \values_reg[12][11]  (.D(values[11]), .CK(n_121_9), .Q(
      \values[12] [11]), .QN());
   DFF_X1 \values_reg[12][10]  (.D(values[10]), .CK(n_121_9), .Q(
      \values[12] [10]), .QN());
   DFF_X1 \values_reg[12][9]  (.D(values[9]), .CK(n_121_9), .Q(\values[12] [9]), 
      .QN());
   DFF_X1 \values_reg[12][8]  (.D(values[8]), .CK(n_121_9), .Q(\values[12] [8]), 
      .QN());
   DFF_X1 \values_reg[12][7]  (.D(values[7]), .CK(n_121_9), .Q(\values[12] [7]), 
      .QN());
   DFF_X1 \values_reg[12][6]  (.D(values[6]), .CK(n_121_9), .Q(\values[12] [6]), 
      .QN());
   DFF_X1 \values_reg[12][5]  (.D(values[5]), .CK(n_121_9), .Q(\values[12] [5]), 
      .QN());
   DFF_X1 \values_reg[12][4]  (.D(values[4]), .CK(n_121_9), .Q(\values[12] [4]), 
      .QN());
   DFF_X1 \values_reg[12][3]  (.D(values[3]), .CK(n_121_9), .Q(\values[12] [3]), 
      .QN());
   DFF_X1 \values_reg[12][2]  (.D(values[2]), .CK(n_121_9), .Q(\values[12] [2]), 
      .QN());
   DFF_X1 \values_reg[12][1]  (.D(values[1]), .CK(n_121_9), .Q(\values[12] [1]), 
      .QN());
   DFF_X1 \values_reg[12][0]  (.D(values[0]), .CK(n_121_9), .Q(\values[12] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[13]_reg  (.CK(clk), .E(n_13), .SE(1'b0), 
      .GCK(n_121_10));
   DFF_X1 \values_reg[13][15]  (.D(values[15]), .CK(n_121_10), .Q(
      \values[13] [15]), .QN());
   DFF_X1 \values_reg[13][14]  (.D(values[14]), .CK(n_121_10), .Q(
      \values[13] [14]), .QN());
   DFF_X1 \values_reg[13][13]  (.D(values[13]), .CK(n_121_10), .Q(
      \values[13] [13]), .QN());
   DFF_X1 \values_reg[13][12]  (.D(values[12]), .CK(n_121_10), .Q(
      \values[13] [12]), .QN());
   DFF_X1 \values_reg[13][11]  (.D(values[11]), .CK(n_121_10), .Q(
      \values[13] [11]), .QN());
   DFF_X1 \values_reg[13][10]  (.D(values[10]), .CK(n_121_10), .Q(
      \values[13] [10]), .QN());
   DFF_X1 \values_reg[13][9]  (.D(values[9]), .CK(n_121_10), .Q(\values[13] [9]), 
      .QN());
   DFF_X1 \values_reg[13][8]  (.D(values[8]), .CK(n_121_10), .Q(\values[13] [8]), 
      .QN());
   DFF_X1 \values_reg[13][7]  (.D(values[7]), .CK(n_121_10), .Q(\values[13] [7]), 
      .QN());
   DFF_X1 \values_reg[13][6]  (.D(values[6]), .CK(n_121_10), .Q(\values[13] [6]), 
      .QN());
   DFF_X1 \values_reg[13][5]  (.D(values[5]), .CK(n_121_10), .Q(\values[13] [5]), 
      .QN());
   DFF_X1 \values_reg[13][4]  (.D(values[4]), .CK(n_121_10), .Q(\values[13] [4]), 
      .QN());
   DFF_X1 \values_reg[13][3]  (.D(values[3]), .CK(n_121_10), .Q(\values[13] [3]), 
      .QN());
   DFF_X1 \values_reg[13][2]  (.D(values[2]), .CK(n_121_10), .Q(\values[13] [2]), 
      .QN());
   DFF_X1 \values_reg[13][1]  (.D(values[1]), .CK(n_121_10), .Q(\values[13] [1]), 
      .QN());
   DFF_X1 \values_reg[13][0]  (.D(values[0]), .CK(n_121_10), .Q(\values[13] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[14]_reg  (.CK(clk), .E(n_14), .SE(1'b0), 
      .GCK(n_121_11));
   DFF_X1 \values_reg[14][15]  (.D(values[15]), .CK(n_121_11), .Q(
      \values[14] [15]), .QN());
   DFF_X1 \values_reg[14][14]  (.D(values[14]), .CK(n_121_11), .Q(
      \values[14] [14]), .QN());
   DFF_X1 \values_reg[14][13]  (.D(values[13]), .CK(n_121_11), .Q(
      \values[14] [13]), .QN());
   DFF_X1 \values_reg[14][12]  (.D(values[12]), .CK(n_121_11), .Q(
      \values[14] [12]), .QN());
   DFF_X1 \values_reg[14][11]  (.D(values[11]), .CK(n_121_11), .Q(
      \values[14] [11]), .QN());
   DFF_X1 \values_reg[14][10]  (.D(values[10]), .CK(n_121_11), .Q(
      \values[14] [10]), .QN());
   DFF_X1 \values_reg[14][9]  (.D(values[9]), .CK(n_121_11), .Q(\values[14] [9]), 
      .QN());
   DFF_X1 \values_reg[14][8]  (.D(values[8]), .CK(n_121_11), .Q(\values[14] [8]), 
      .QN());
   DFF_X1 \values_reg[14][7]  (.D(values[7]), .CK(n_121_11), .Q(\values[14] [7]), 
      .QN());
   DFF_X1 \values_reg[14][6]  (.D(values[6]), .CK(n_121_11), .Q(\values[14] [6]), 
      .QN());
   DFF_X1 \values_reg[14][5]  (.D(values[5]), .CK(n_121_11), .Q(\values[14] [5]), 
      .QN());
   DFF_X1 \values_reg[14][4]  (.D(values[4]), .CK(n_121_11), .Q(\values[14] [4]), 
      .QN());
   DFF_X1 \values_reg[14][3]  (.D(values[3]), .CK(n_121_11), .Q(\values[14] [3]), 
      .QN());
   DFF_X1 \values_reg[14][2]  (.D(values[2]), .CK(n_121_11), .Q(\values[14] [2]), 
      .QN());
   DFF_X1 \values_reg[14][1]  (.D(values[1]), .CK(n_121_11), .Q(\values[14] [1]), 
      .QN());
   DFF_X1 \values_reg[14][0]  (.D(values[0]), .CK(n_121_11), .Q(\values[14] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[15]_reg  (.CK(clk), .E(n_15), .SE(1'b0), 
      .GCK(n_121_12));
   DFF_X1 \values_reg[15][15]  (.D(values[15]), .CK(n_121_12), .Q(
      \values[15] [15]), .QN());
   DFF_X1 \values_reg[15][14]  (.D(values[14]), .CK(n_121_12), .Q(
      \values[15] [14]), .QN());
   DFF_X1 \values_reg[15][13]  (.D(values[13]), .CK(n_121_12), .Q(
      \values[15] [13]), .QN());
   DFF_X1 \values_reg[15][12]  (.D(values[12]), .CK(n_121_12), .Q(
      \values[15] [12]), .QN());
   DFF_X1 \values_reg[15][11]  (.D(values[11]), .CK(n_121_12), .Q(
      \values[15] [11]), .QN());
   DFF_X1 \values_reg[15][10]  (.D(values[10]), .CK(n_121_12), .Q(
      \values[15] [10]), .QN());
   DFF_X1 \values_reg[15][9]  (.D(values[9]), .CK(n_121_12), .Q(\values[15] [9]), 
      .QN());
   DFF_X1 \values_reg[15][8]  (.D(values[8]), .CK(n_121_12), .Q(\values[15] [8]), 
      .QN());
   DFF_X1 \values_reg[15][7]  (.D(values[7]), .CK(n_121_12), .Q(\values[15] [7]), 
      .QN());
   DFF_X1 \values_reg[15][6]  (.D(values[6]), .CK(n_121_12), .Q(\values[15] [6]), 
      .QN());
   DFF_X1 \values_reg[15][5]  (.D(values[5]), .CK(n_121_12), .Q(\values[15] [5]), 
      .QN());
   DFF_X1 \values_reg[15][4]  (.D(values[4]), .CK(n_121_12), .Q(\values[15] [4]), 
      .QN());
   DFF_X1 \values_reg[15][3]  (.D(values[3]), .CK(n_121_12), .Q(\values[15] [3]), 
      .QN());
   DFF_X1 \values_reg[15][2]  (.D(values[2]), .CK(n_121_12), .Q(\values[15] [2]), 
      .QN());
   DFF_X1 \values_reg[15][1]  (.D(values[1]), .CK(n_121_12), .Q(\values[15] [1]), 
      .QN());
   DFF_X1 \values_reg[15][0]  (.D(values[0]), .CK(n_121_12), .Q(\values[15] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[16]_reg  (.CK(clk), .E(n_16), .SE(1'b0), 
      .GCK(n_121_13));
   DFF_X1 \values_reg[16][15]  (.D(values[15]), .CK(n_121_13), .Q(
      \values[16] [15]), .QN());
   DFF_X1 \values_reg[16][14]  (.D(values[14]), .CK(n_121_13), .Q(
      \values[16] [14]), .QN());
   DFF_X1 \values_reg[16][13]  (.D(values[13]), .CK(n_121_13), .Q(
      \values[16] [13]), .QN());
   DFF_X1 \values_reg[16][12]  (.D(values[12]), .CK(n_121_13), .Q(
      \values[16] [12]), .QN());
   DFF_X1 \values_reg[16][11]  (.D(values[11]), .CK(n_121_13), .Q(
      \values[16] [11]), .QN());
   DFF_X1 \values_reg[16][10]  (.D(values[10]), .CK(n_121_13), .Q(
      \values[16] [10]), .QN());
   DFF_X1 \values_reg[16][9]  (.D(values[9]), .CK(n_121_13), .Q(\values[16] [9]), 
      .QN());
   DFF_X1 \values_reg[16][8]  (.D(values[8]), .CK(n_121_13), .Q(\values[16] [8]), 
      .QN());
   DFF_X1 \values_reg[16][7]  (.D(values[7]), .CK(n_121_13), .Q(\values[16] [7]), 
      .QN());
   DFF_X1 \values_reg[16][6]  (.D(values[6]), .CK(n_121_13), .Q(\values[16] [6]), 
      .QN());
   DFF_X1 \values_reg[16][5]  (.D(values[5]), .CK(n_121_13), .Q(\values[16] [5]), 
      .QN());
   DFF_X1 \values_reg[16][4]  (.D(values[4]), .CK(n_121_13), .Q(\values[16] [4]), 
      .QN());
   DFF_X1 \values_reg[16][3]  (.D(values[3]), .CK(n_121_13), .Q(\values[16] [3]), 
      .QN());
   DFF_X1 \values_reg[16][2]  (.D(values[2]), .CK(n_121_13), .Q(\values[16] [2]), 
      .QN());
   DFF_X1 \values_reg[16][1]  (.D(values[1]), .CK(n_121_13), .Q(\values[16] [1]), 
      .QN());
   DFF_X1 \values_reg[16][0]  (.D(values[0]), .CK(n_121_13), .Q(\values[16] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[17]_reg  (.CK(clk), .E(n_17), .SE(1'b0), 
      .GCK(n_121_14));
   DFF_X1 \values_reg[17][15]  (.D(values[15]), .CK(n_121_14), .Q(
      \values[17] [15]), .QN());
   DFF_X1 \values_reg[17][14]  (.D(values[14]), .CK(n_121_14), .Q(
      \values[17] [14]), .QN());
   DFF_X1 \values_reg[17][13]  (.D(values[13]), .CK(n_121_14), .Q(
      \values[17] [13]), .QN());
   DFF_X1 \values_reg[17][12]  (.D(values[12]), .CK(n_121_14), .Q(
      \values[17] [12]), .QN());
   DFF_X1 \values_reg[17][11]  (.D(values[11]), .CK(n_121_14), .Q(
      \values[17] [11]), .QN());
   DFF_X1 \values_reg[17][10]  (.D(values[10]), .CK(n_121_14), .Q(
      \values[17] [10]), .QN());
   DFF_X1 \values_reg[17][9]  (.D(values[9]), .CK(n_121_14), .Q(\values[17] [9]), 
      .QN());
   DFF_X1 \values_reg[17][8]  (.D(values[8]), .CK(n_121_14), .Q(\values[17] [8]), 
      .QN());
   DFF_X1 \values_reg[17][7]  (.D(values[7]), .CK(n_121_14), .Q(\values[17] [7]), 
      .QN());
   DFF_X1 \values_reg[17][6]  (.D(values[6]), .CK(n_121_14), .Q(\values[17] [6]), 
      .QN());
   DFF_X1 \values_reg[17][5]  (.D(values[5]), .CK(n_121_14), .Q(\values[17] [5]), 
      .QN());
   DFF_X1 \values_reg[17][4]  (.D(values[4]), .CK(n_121_14), .Q(\values[17] [4]), 
      .QN());
   DFF_X1 \values_reg[17][3]  (.D(values[3]), .CK(n_121_14), .Q(\values[17] [3]), 
      .QN());
   DFF_X1 \values_reg[17][2]  (.D(values[2]), .CK(n_121_14), .Q(\values[17] [2]), 
      .QN());
   DFF_X1 \values_reg[17][1]  (.D(values[1]), .CK(n_121_14), .Q(\values[17] [1]), 
      .QN());
   DFF_X1 \values_reg[17][0]  (.D(values[0]), .CK(n_121_14), .Q(\values[17] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[18]_reg  (.CK(clk), .E(n_18), .SE(1'b0), 
      .GCK(n_121_15));
   DFF_X1 \values_reg[18][15]  (.D(values[15]), .CK(n_121_15), .Q(
      \values[18] [15]), .QN());
   DFF_X1 \values_reg[18][14]  (.D(values[14]), .CK(n_121_15), .Q(
      \values[18] [14]), .QN());
   DFF_X1 \values_reg[18][13]  (.D(values[13]), .CK(n_121_15), .Q(
      \values[18] [13]), .QN());
   DFF_X1 \values_reg[18][12]  (.D(values[12]), .CK(n_121_15), .Q(
      \values[18] [12]), .QN());
   DFF_X1 \values_reg[18][11]  (.D(values[11]), .CK(n_121_15), .Q(
      \values[18] [11]), .QN());
   DFF_X1 \values_reg[18][10]  (.D(values[10]), .CK(n_121_15), .Q(
      \values[18] [10]), .QN());
   DFF_X1 \values_reg[18][9]  (.D(values[9]), .CK(n_121_15), .Q(\values[18] [9]), 
      .QN());
   DFF_X1 \values_reg[18][8]  (.D(values[8]), .CK(n_121_15), .Q(\values[18] [8]), 
      .QN());
   DFF_X1 \values_reg[18][7]  (.D(values[7]), .CK(n_121_15), .Q(\values[18] [7]), 
      .QN());
   DFF_X1 \values_reg[18][6]  (.D(values[6]), .CK(n_121_15), .Q(\values[18] [6]), 
      .QN());
   DFF_X1 \values_reg[18][5]  (.D(values[5]), .CK(n_121_15), .Q(\values[18] [5]), 
      .QN());
   DFF_X1 \values_reg[18][4]  (.D(values[4]), .CK(n_121_15), .Q(\values[18] [4]), 
      .QN());
   DFF_X1 \values_reg[18][3]  (.D(values[3]), .CK(n_121_15), .Q(\values[18] [3]), 
      .QN());
   DFF_X1 \values_reg[18][2]  (.D(values[2]), .CK(n_121_15), .Q(\values[18] [2]), 
      .QN());
   DFF_X1 \values_reg[18][1]  (.D(values[1]), .CK(n_121_15), .Q(\values[18] [1]), 
      .QN());
   DFF_X1 \values_reg[18][0]  (.D(values[0]), .CK(n_121_15), .Q(\values[18] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[19]_reg  (.CK(clk), .E(n_19), .SE(1'b0), 
      .GCK(n_121_16));
   DFF_X1 \values_reg[19][15]  (.D(values[15]), .CK(n_121_16), .Q(
      \values[19] [15]), .QN());
   DFF_X1 \values_reg[19][14]  (.D(values[14]), .CK(n_121_16), .Q(
      \values[19] [14]), .QN());
   DFF_X1 \values_reg[19][13]  (.D(values[13]), .CK(n_121_16), .Q(
      \values[19] [13]), .QN());
   DFF_X1 \values_reg[19][12]  (.D(values[12]), .CK(n_121_16), .Q(
      \values[19] [12]), .QN());
   DFF_X1 \values_reg[19][11]  (.D(values[11]), .CK(n_121_16), .Q(
      \values[19] [11]), .QN());
   DFF_X1 \values_reg[19][10]  (.D(values[10]), .CK(n_121_16), .Q(
      \values[19] [10]), .QN());
   DFF_X1 \values_reg[19][9]  (.D(values[9]), .CK(n_121_16), .Q(\values[19] [9]), 
      .QN());
   DFF_X1 \values_reg[19][8]  (.D(values[8]), .CK(n_121_16), .Q(\values[19] [8]), 
      .QN());
   DFF_X1 \values_reg[19][7]  (.D(values[7]), .CK(n_121_16), .Q(\values[19] [7]), 
      .QN());
   DFF_X1 \values_reg[19][6]  (.D(values[6]), .CK(n_121_16), .Q(\values[19] [6]), 
      .QN());
   DFF_X1 \values_reg[19][5]  (.D(values[5]), .CK(n_121_16), .Q(\values[19] [5]), 
      .QN());
   DFF_X1 \values_reg[19][4]  (.D(values[4]), .CK(n_121_16), .Q(\values[19] [4]), 
      .QN());
   DFF_X1 \values_reg[19][3]  (.D(values[3]), .CK(n_121_16), .Q(\values[19] [3]), 
      .QN());
   DFF_X1 \values_reg[19][2]  (.D(values[2]), .CK(n_121_16), .Q(\values[19] [2]), 
      .QN());
   DFF_X1 \values_reg[19][1]  (.D(values[1]), .CK(n_121_16), .Q(\values[19] [1]), 
      .QN());
   DFF_X1 \values_reg[19][0]  (.D(values[0]), .CK(n_121_16), .Q(\values[19] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[20]_reg  (.CK(clk), .E(n_20), .SE(1'b0), 
      .GCK(n_121_17));
   DFF_X1 \values_reg[20][15]  (.D(values[15]), .CK(n_121_17), .Q(
      \values[20] [15]), .QN());
   DFF_X1 \values_reg[20][14]  (.D(values[14]), .CK(n_121_17), .Q(
      \values[20] [14]), .QN());
   DFF_X1 \values_reg[20][13]  (.D(values[13]), .CK(n_121_17), .Q(
      \values[20] [13]), .QN());
   DFF_X1 \values_reg[20][12]  (.D(values[12]), .CK(n_121_17), .Q(
      \values[20] [12]), .QN());
   DFF_X1 \values_reg[20][11]  (.D(values[11]), .CK(n_121_17), .Q(
      \values[20] [11]), .QN());
   DFF_X1 \values_reg[20][10]  (.D(values[10]), .CK(n_121_17), .Q(
      \values[20] [10]), .QN());
   DFF_X1 \values_reg[20][9]  (.D(values[9]), .CK(n_121_17), .Q(\values[20] [9]), 
      .QN());
   DFF_X1 \values_reg[20][8]  (.D(values[8]), .CK(n_121_17), .Q(\values[20] [8]), 
      .QN());
   DFF_X1 \values_reg[20][7]  (.D(values[7]), .CK(n_121_17), .Q(\values[20] [7]), 
      .QN());
   DFF_X1 \values_reg[20][6]  (.D(values[6]), .CK(n_121_17), .Q(\values[20] [6]), 
      .QN());
   DFF_X1 \values_reg[20][5]  (.D(values[5]), .CK(n_121_17), .Q(\values[20] [5]), 
      .QN());
   DFF_X1 \values_reg[20][4]  (.D(values[4]), .CK(n_121_17), .Q(\values[20] [4]), 
      .QN());
   DFF_X1 \values_reg[20][3]  (.D(values[3]), .CK(n_121_17), .Q(\values[20] [3]), 
      .QN());
   DFF_X1 \values_reg[20][2]  (.D(values[2]), .CK(n_121_17), .Q(\values[20] [2]), 
      .QN());
   DFF_X1 \values_reg[20][1]  (.D(values[1]), .CK(n_121_17), .Q(\values[20] [1]), 
      .QN());
   DFF_X1 \values_reg[20][0]  (.D(values[0]), .CK(n_121_17), .Q(\values[20] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[21]_reg  (.CK(clk), .E(n_21), .SE(1'b0), 
      .GCK(n_121_18));
   DFF_X1 \values_reg[21][15]  (.D(values[15]), .CK(n_121_18), .Q(
      \values[21] [15]), .QN());
   DFF_X1 \values_reg[21][14]  (.D(values[14]), .CK(n_121_18), .Q(
      \values[21] [14]), .QN());
   DFF_X1 \values_reg[21][13]  (.D(values[13]), .CK(n_121_18), .Q(
      \values[21] [13]), .QN());
   DFF_X1 \values_reg[21][12]  (.D(values[12]), .CK(n_121_18), .Q(
      \values[21] [12]), .QN());
   DFF_X1 \values_reg[21][11]  (.D(values[11]), .CK(n_121_18), .Q(
      \values[21] [11]), .QN());
   DFF_X1 \values_reg[21][10]  (.D(values[10]), .CK(n_121_18), .Q(
      \values[21] [10]), .QN());
   DFF_X1 \values_reg[21][9]  (.D(values[9]), .CK(n_121_18), .Q(\values[21] [9]), 
      .QN());
   DFF_X1 \values_reg[21][8]  (.D(values[8]), .CK(n_121_18), .Q(\values[21] [8]), 
      .QN());
   DFF_X1 \values_reg[21][7]  (.D(values[7]), .CK(n_121_18), .Q(\values[21] [7]), 
      .QN());
   DFF_X1 \values_reg[21][6]  (.D(values[6]), .CK(n_121_18), .Q(\values[21] [6]), 
      .QN());
   DFF_X1 \values_reg[21][5]  (.D(values[5]), .CK(n_121_18), .Q(\values[21] [5]), 
      .QN());
   DFF_X1 \values_reg[21][4]  (.D(values[4]), .CK(n_121_18), .Q(\values[21] [4]), 
      .QN());
   DFF_X1 \values_reg[21][3]  (.D(values[3]), .CK(n_121_18), .Q(\values[21] [3]), 
      .QN());
   DFF_X1 \values_reg[21][2]  (.D(values[2]), .CK(n_121_18), .Q(\values[21] [2]), 
      .QN());
   DFF_X1 \values_reg[21][1]  (.D(values[1]), .CK(n_121_18), .Q(\values[21] [1]), 
      .QN());
   DFF_X1 \values_reg[21][0]  (.D(values[0]), .CK(n_121_18), .Q(\values[21] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[22]_reg  (.CK(clk), .E(n_22), .SE(1'b0), 
      .GCK(n_121_19));
   DFF_X1 \values_reg[22][15]  (.D(values[15]), .CK(n_121_19), .Q(
      \values[22] [15]), .QN());
   DFF_X1 \values_reg[22][14]  (.D(values[14]), .CK(n_121_19), .Q(
      \values[22] [14]), .QN());
   DFF_X1 \values_reg[22][13]  (.D(values[13]), .CK(n_121_19), .Q(
      \values[22] [13]), .QN());
   DFF_X1 \values_reg[22][12]  (.D(values[12]), .CK(n_121_19), .Q(
      \values[22] [12]), .QN());
   DFF_X1 \values_reg[22][11]  (.D(values[11]), .CK(n_121_19), .Q(
      \values[22] [11]), .QN());
   DFF_X1 \values_reg[22][10]  (.D(values[10]), .CK(n_121_19), .Q(
      \values[22] [10]), .QN());
   DFF_X1 \values_reg[22][9]  (.D(values[9]), .CK(n_121_19), .Q(\values[22] [9]), 
      .QN());
   DFF_X1 \values_reg[22][8]  (.D(values[8]), .CK(n_121_19), .Q(\values[22] [8]), 
      .QN());
   DFF_X1 \values_reg[22][7]  (.D(values[7]), .CK(n_121_19), .Q(\values[22] [7]), 
      .QN());
   DFF_X1 \values_reg[22][6]  (.D(values[6]), .CK(n_121_19), .Q(\values[22] [6]), 
      .QN());
   DFF_X1 \values_reg[22][5]  (.D(values[5]), .CK(n_121_19), .Q(\values[22] [5]), 
      .QN());
   DFF_X1 \values_reg[22][4]  (.D(values[4]), .CK(n_121_19), .Q(\values[22] [4]), 
      .QN());
   DFF_X1 \values_reg[22][3]  (.D(values[3]), .CK(n_121_19), .Q(\values[22] [3]), 
      .QN());
   DFF_X1 \values_reg[22][2]  (.D(values[2]), .CK(n_121_19), .Q(\values[22] [2]), 
      .QN());
   DFF_X1 \values_reg[22][1]  (.D(values[1]), .CK(n_121_19), .Q(\values[22] [1]), 
      .QN());
   DFF_X1 \values_reg[22][0]  (.D(values[0]), .CK(n_121_19), .Q(\values[22] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[23]_reg  (.CK(clk), .E(n_23), .SE(1'b0), 
      .GCK(n_121_20));
   DFF_X1 \values_reg[23][15]  (.D(values[15]), .CK(n_121_20), .Q(
      \values[23] [15]), .QN());
   DFF_X1 \values_reg[23][14]  (.D(values[14]), .CK(n_121_20), .Q(
      \values[23] [14]), .QN());
   DFF_X1 \values_reg[23][13]  (.D(values[13]), .CK(n_121_20), .Q(
      \values[23] [13]), .QN());
   DFF_X1 \values_reg[23][12]  (.D(values[12]), .CK(n_121_20), .Q(
      \values[23] [12]), .QN());
   DFF_X1 \values_reg[23][11]  (.D(values[11]), .CK(n_121_20), .Q(
      \values[23] [11]), .QN());
   DFF_X1 \values_reg[23][10]  (.D(values[10]), .CK(n_121_20), .Q(
      \values[23] [10]), .QN());
   DFF_X1 \values_reg[23][9]  (.D(values[9]), .CK(n_121_20), .Q(\values[23] [9]), 
      .QN());
   DFF_X1 \values_reg[23][8]  (.D(values[8]), .CK(n_121_20), .Q(\values[23] [8]), 
      .QN());
   DFF_X1 \values_reg[23][7]  (.D(values[7]), .CK(n_121_20), .Q(\values[23] [7]), 
      .QN());
   DFF_X1 \values_reg[23][6]  (.D(values[6]), .CK(n_121_20), .Q(\values[23] [6]), 
      .QN());
   DFF_X1 \values_reg[23][5]  (.D(values[5]), .CK(n_121_20), .Q(\values[23] [5]), 
      .QN());
   DFF_X1 \values_reg[23][4]  (.D(values[4]), .CK(n_121_20), .Q(\values[23] [4]), 
      .QN());
   DFF_X1 \values_reg[23][3]  (.D(values[3]), .CK(n_121_20), .Q(\values[23] [3]), 
      .QN());
   DFF_X1 \values_reg[23][2]  (.D(values[2]), .CK(n_121_20), .Q(\values[23] [2]), 
      .QN());
   DFF_X1 \values_reg[23][1]  (.D(values[1]), .CK(n_121_20), .Q(\values[23] [1]), 
      .QN());
   DFF_X1 \values_reg[23][0]  (.D(values[0]), .CK(n_121_20), .Q(\values[23] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[24]_reg  (.CK(clk), .E(n_24), .SE(1'b0), 
      .GCK(n_121_21));
   DFF_X1 \values_reg[24][15]  (.D(values[15]), .CK(n_121_21), .Q(
      \values[24] [15]), .QN());
   DFF_X1 \values_reg[24][14]  (.D(values[14]), .CK(n_121_21), .Q(
      \values[24] [14]), .QN());
   DFF_X1 \values_reg[24][13]  (.D(values[13]), .CK(n_121_21), .Q(
      \values[24] [13]), .QN());
   DFF_X1 \values_reg[24][12]  (.D(values[12]), .CK(n_121_21), .Q(
      \values[24] [12]), .QN());
   DFF_X1 \values_reg[24][11]  (.D(values[11]), .CK(n_121_21), .Q(
      \values[24] [11]), .QN());
   DFF_X1 \values_reg[24][10]  (.D(values[10]), .CK(n_121_21), .Q(
      \values[24] [10]), .QN());
   DFF_X1 \values_reg[24][9]  (.D(values[9]), .CK(n_121_21), .Q(\values[24] [9]), 
      .QN());
   DFF_X1 \values_reg[24][8]  (.D(values[8]), .CK(n_121_21), .Q(\values[24] [8]), 
      .QN());
   DFF_X1 \values_reg[24][7]  (.D(values[7]), .CK(n_121_21), .Q(\values[24] [7]), 
      .QN());
   DFF_X1 \values_reg[24][6]  (.D(values[6]), .CK(n_121_21), .Q(\values[24] [6]), 
      .QN());
   DFF_X1 \values_reg[24][5]  (.D(values[5]), .CK(n_121_21), .Q(\values[24] [5]), 
      .QN());
   DFF_X1 \values_reg[24][4]  (.D(values[4]), .CK(n_121_21), .Q(\values[24] [4]), 
      .QN());
   DFF_X1 \values_reg[24][3]  (.D(values[3]), .CK(n_121_21), .Q(\values[24] [3]), 
      .QN());
   DFF_X1 \values_reg[24][2]  (.D(values[2]), .CK(n_121_21), .Q(\values[24] [2]), 
      .QN());
   DFF_X1 \values_reg[24][1]  (.D(values[1]), .CK(n_121_21), .Q(\values[24] [1]), 
      .QN());
   DFF_X1 \values_reg[24][0]  (.D(values[0]), .CK(n_121_21), .Q(\values[24] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[25]_reg  (.CK(clk), .E(n_25), .SE(1'b0), 
      .GCK(n_121_22));
   DFF_X1 \values_reg[25][15]  (.D(values[15]), .CK(n_121_22), .Q(
      \values[25] [15]), .QN());
   DFF_X1 \values_reg[25][14]  (.D(values[14]), .CK(n_121_22), .Q(
      \values[25] [14]), .QN());
   DFF_X1 \values_reg[25][13]  (.D(values[13]), .CK(n_121_22), .Q(
      \values[25] [13]), .QN());
   DFF_X1 \values_reg[25][12]  (.D(values[12]), .CK(n_121_22), .Q(
      \values[25] [12]), .QN());
   DFF_X1 \values_reg[25][11]  (.D(values[11]), .CK(n_121_22), .Q(
      \values[25] [11]), .QN());
   DFF_X1 \values_reg[25][10]  (.D(values[10]), .CK(n_121_22), .Q(
      \values[25] [10]), .QN());
   DFF_X1 \values_reg[25][9]  (.D(values[9]), .CK(n_121_22), .Q(\values[25] [9]), 
      .QN());
   DFF_X1 \values_reg[25][8]  (.D(values[8]), .CK(n_121_22), .Q(\values[25] [8]), 
      .QN());
   DFF_X1 \values_reg[25][7]  (.D(values[7]), .CK(n_121_22), .Q(\values[25] [7]), 
      .QN());
   DFF_X1 \values_reg[25][6]  (.D(values[6]), .CK(n_121_22), .Q(\values[25] [6]), 
      .QN());
   DFF_X1 \values_reg[25][5]  (.D(values[5]), .CK(n_121_22), .Q(\values[25] [5]), 
      .QN());
   DFF_X1 \values_reg[25][4]  (.D(values[4]), .CK(n_121_22), .Q(\values[25] [4]), 
      .QN());
   DFF_X1 \values_reg[25][3]  (.D(values[3]), .CK(n_121_22), .Q(\values[25] [3]), 
      .QN());
   DFF_X1 \values_reg[25][2]  (.D(values[2]), .CK(n_121_22), .Q(\values[25] [2]), 
      .QN());
   DFF_X1 \values_reg[25][1]  (.D(values[1]), .CK(n_121_22), .Q(\values[25] [1]), 
      .QN());
   DFF_X1 \values_reg[25][0]  (.D(values[0]), .CK(n_121_22), .Q(\values[25] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[96]_reg  (.CK(clk), .E(n_96), .SE(1'b0), 
      .GCK(n_121_23));
   DFF_X1 \values_reg[96][15]  (.D(values[15]), .CK(n_121_23), .Q(
      \values[96] [15]), .QN());
   DFF_X1 \values_reg[96][14]  (.D(values[14]), .CK(n_121_23), .Q(
      \values[96] [14]), .QN());
   DFF_X1 \values_reg[96][13]  (.D(values[13]), .CK(n_121_23), .Q(
      \values[96] [13]), .QN());
   DFF_X1 \values_reg[96][12]  (.D(values[12]), .CK(n_121_23), .Q(
      \values[96] [12]), .QN());
   DFF_X1 \values_reg[96][11]  (.D(values[11]), .CK(n_121_23), .Q(
      \values[96] [11]), .QN());
   DFF_X1 \values_reg[96][10]  (.D(values[10]), .CK(n_121_23), .Q(
      \values[96] [10]), .QN());
   DFF_X1 \values_reg[96][9]  (.D(values[9]), .CK(n_121_23), .Q(\values[96] [9]), 
      .QN());
   DFF_X1 \values_reg[96][8]  (.D(values[8]), .CK(n_121_23), .Q(\values[96] [8]), 
      .QN());
   DFF_X1 \values_reg[96][7]  (.D(values[7]), .CK(n_121_23), .Q(\values[96] [7]), 
      .QN());
   DFF_X1 \values_reg[96][6]  (.D(values[6]), .CK(n_121_23), .Q(\values[96] [6]), 
      .QN());
   DFF_X1 \values_reg[96][5]  (.D(values[5]), .CK(n_121_23), .Q(\values[96] [5]), 
      .QN());
   DFF_X1 \values_reg[96][4]  (.D(values[4]), .CK(n_121_23), .Q(\values[96] [4]), 
      .QN());
   DFF_X1 \values_reg[96][3]  (.D(values[3]), .CK(n_121_23), .Q(\values[96] [3]), 
      .QN());
   DFF_X1 \values_reg[96][2]  (.D(values[2]), .CK(n_121_23), .Q(\values[96] [2]), 
      .QN());
   DFF_X1 \values_reg[96][1]  (.D(values[1]), .CK(n_121_23), .Q(\values[96] [1]), 
      .QN());
   DFF_X1 \values_reg[96][0]  (.D(values[0]), .CK(n_121_23), .Q(\values[96] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[95]_reg  (.CK(clk), .E(n_95), .SE(1'b0), 
      .GCK(n_121_24));
   DFF_X1 \values_reg[95][15]  (.D(values[15]), .CK(n_121_24), .Q(
      \values[95] [15]), .QN());
   DFF_X1 \values_reg[95][14]  (.D(values[14]), .CK(n_121_24), .Q(
      \values[95] [14]), .QN());
   DFF_X1 \values_reg[95][13]  (.D(values[13]), .CK(n_121_24), .Q(
      \values[95] [13]), .QN());
   DFF_X1 \values_reg[95][12]  (.D(values[12]), .CK(n_121_24), .Q(
      \values[95] [12]), .QN());
   DFF_X1 \values_reg[95][11]  (.D(values[11]), .CK(n_121_24), .Q(
      \values[95] [11]), .QN());
   DFF_X1 \values_reg[95][10]  (.D(values[10]), .CK(n_121_24), .Q(
      \values[95] [10]), .QN());
   DFF_X1 \values_reg[95][9]  (.D(values[9]), .CK(n_121_24), .Q(\values[95] [9]), 
      .QN());
   DFF_X1 \values_reg[95][8]  (.D(values[8]), .CK(n_121_24), .Q(\values[95] [8]), 
      .QN());
   DFF_X1 \values_reg[95][7]  (.D(values[7]), .CK(n_121_24), .Q(\values[95] [7]), 
      .QN());
   DFF_X1 \values_reg[95][6]  (.D(values[6]), .CK(n_121_24), .Q(\values[95] [6]), 
      .QN());
   DFF_X1 \values_reg[95][5]  (.D(values[5]), .CK(n_121_24), .Q(\values[95] [5]), 
      .QN());
   DFF_X1 \values_reg[95][4]  (.D(values[4]), .CK(n_121_24), .Q(\values[95] [4]), 
      .QN());
   DFF_X1 \values_reg[95][3]  (.D(values[3]), .CK(n_121_24), .Q(\values[95] [3]), 
      .QN());
   DFF_X1 \values_reg[95][2]  (.D(values[2]), .CK(n_121_24), .Q(\values[95] [2]), 
      .QN());
   DFF_X1 \values_reg[95][1]  (.D(values[1]), .CK(n_121_24), .Q(\values[95] [1]), 
      .QN());
   DFF_X1 \values_reg[95][0]  (.D(values[0]), .CK(n_121_24), .Q(\values[95] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[94]_reg  (.CK(clk), .E(n_94), .SE(1'b0), 
      .GCK(n_121_25));
   DFF_X1 \values_reg[94][15]  (.D(values[15]), .CK(n_121_25), .Q(
      \values[94] [15]), .QN());
   DFF_X1 \values_reg[94][14]  (.D(values[14]), .CK(n_121_25), .Q(
      \values[94] [14]), .QN());
   DFF_X1 \values_reg[94][13]  (.D(values[13]), .CK(n_121_25), .Q(
      \values[94] [13]), .QN());
   DFF_X1 \values_reg[94][12]  (.D(values[12]), .CK(n_121_25), .Q(
      \values[94] [12]), .QN());
   DFF_X1 \values_reg[94][11]  (.D(values[11]), .CK(n_121_25), .Q(
      \values[94] [11]), .QN());
   DFF_X1 \values_reg[94][10]  (.D(values[10]), .CK(n_121_25), .Q(
      \values[94] [10]), .QN());
   DFF_X1 \values_reg[94][9]  (.D(values[9]), .CK(n_121_25), .Q(\values[94] [9]), 
      .QN());
   DFF_X1 \values_reg[94][8]  (.D(values[8]), .CK(n_121_25), .Q(\values[94] [8]), 
      .QN());
   DFF_X1 \values_reg[94][7]  (.D(values[7]), .CK(n_121_25), .Q(\values[94] [7]), 
      .QN());
   DFF_X1 \values_reg[94][6]  (.D(values[6]), .CK(n_121_25), .Q(\values[94] [6]), 
      .QN());
   DFF_X1 \values_reg[94][5]  (.D(values[5]), .CK(n_121_25), .Q(\values[94] [5]), 
      .QN());
   DFF_X1 \values_reg[94][4]  (.D(values[4]), .CK(n_121_25), .Q(\values[94] [4]), 
      .QN());
   DFF_X1 \values_reg[94][3]  (.D(values[3]), .CK(n_121_25), .Q(\values[94] [3]), 
      .QN());
   DFF_X1 \values_reg[94][2]  (.D(values[2]), .CK(n_121_25), .Q(\values[94] [2]), 
      .QN());
   DFF_X1 \values_reg[94][1]  (.D(values[1]), .CK(n_121_25), .Q(\values[94] [1]), 
      .QN());
   DFF_X1 \values_reg[94][0]  (.D(values[0]), .CK(n_121_25), .Q(\values[94] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[93]_reg  (.CK(clk), .E(n_93), .SE(1'b0), 
      .GCK(n_121_26));
   DFF_X1 \values_reg[93][15]  (.D(values[15]), .CK(n_121_26), .Q(
      \values[93] [15]), .QN());
   DFF_X1 \values_reg[93][14]  (.D(values[14]), .CK(n_121_26), .Q(
      \values[93] [14]), .QN());
   DFF_X1 \values_reg[93][13]  (.D(values[13]), .CK(n_121_26), .Q(
      \values[93] [13]), .QN());
   DFF_X1 \values_reg[93][12]  (.D(values[12]), .CK(n_121_26), .Q(
      \values[93] [12]), .QN());
   DFF_X1 \values_reg[93][11]  (.D(values[11]), .CK(n_121_26), .Q(
      \values[93] [11]), .QN());
   DFF_X1 \values_reg[93][10]  (.D(values[10]), .CK(n_121_26), .Q(
      \values[93] [10]), .QN());
   DFF_X1 \values_reg[93][9]  (.D(values[9]), .CK(n_121_26), .Q(\values[93] [9]), 
      .QN());
   DFF_X1 \values_reg[93][8]  (.D(values[8]), .CK(n_121_26), .Q(\values[93] [8]), 
      .QN());
   DFF_X1 \values_reg[93][7]  (.D(values[7]), .CK(n_121_26), .Q(\values[93] [7]), 
      .QN());
   DFF_X1 \values_reg[93][6]  (.D(values[6]), .CK(n_121_26), .Q(\values[93] [6]), 
      .QN());
   DFF_X1 \values_reg[93][5]  (.D(values[5]), .CK(n_121_26), .Q(\values[93] [5]), 
      .QN());
   DFF_X1 \values_reg[93][4]  (.D(values[4]), .CK(n_121_26), .Q(\values[93] [4]), 
      .QN());
   DFF_X1 \values_reg[93][3]  (.D(values[3]), .CK(n_121_26), .Q(\values[93] [3]), 
      .QN());
   DFF_X1 \values_reg[93][2]  (.D(values[2]), .CK(n_121_26), .Q(\values[93] [2]), 
      .QN());
   DFF_X1 \values_reg[93][1]  (.D(values[1]), .CK(n_121_26), .Q(\values[93] [1]), 
      .QN());
   DFF_X1 \values_reg[93][0]  (.D(values[0]), .CK(n_121_26), .Q(\values[93] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[92]_reg  (.CK(clk), .E(n_92), .SE(1'b0), 
      .GCK(n_121_27));
   DFF_X1 \values_reg[92][15]  (.D(values[15]), .CK(n_121_27), .Q(
      \values[92] [15]), .QN());
   DFF_X1 \values_reg[92][14]  (.D(values[14]), .CK(n_121_27), .Q(
      \values[92] [14]), .QN());
   DFF_X1 \values_reg[92][13]  (.D(values[13]), .CK(n_121_27), .Q(
      \values[92] [13]), .QN());
   DFF_X1 \values_reg[92][12]  (.D(values[12]), .CK(n_121_27), .Q(
      \values[92] [12]), .QN());
   DFF_X1 \values_reg[92][11]  (.D(values[11]), .CK(n_121_27), .Q(
      \values[92] [11]), .QN());
   DFF_X1 \values_reg[92][10]  (.D(values[10]), .CK(n_121_27), .Q(
      \values[92] [10]), .QN());
   DFF_X1 \values_reg[92][9]  (.D(values[9]), .CK(n_121_27), .Q(\values[92] [9]), 
      .QN());
   DFF_X1 \values_reg[92][8]  (.D(values[8]), .CK(n_121_27), .Q(\values[92] [8]), 
      .QN());
   DFF_X1 \values_reg[92][7]  (.D(values[7]), .CK(n_121_27), .Q(\values[92] [7]), 
      .QN());
   DFF_X1 \values_reg[92][6]  (.D(values[6]), .CK(n_121_27), .Q(\values[92] [6]), 
      .QN());
   DFF_X1 \values_reg[92][5]  (.D(values[5]), .CK(n_121_27), .Q(\values[92] [5]), 
      .QN());
   DFF_X1 \values_reg[92][4]  (.D(values[4]), .CK(n_121_27), .Q(\values[92] [4]), 
      .QN());
   DFF_X1 \values_reg[92][3]  (.D(values[3]), .CK(n_121_27), .Q(\values[92] [3]), 
      .QN());
   DFF_X1 \values_reg[92][2]  (.D(values[2]), .CK(n_121_27), .Q(\values[92] [2]), 
      .QN());
   DFF_X1 \values_reg[92][1]  (.D(values[1]), .CK(n_121_27), .Q(\values[92] [1]), 
      .QN());
   DFF_X1 \values_reg[92][0]  (.D(values[0]), .CK(n_121_27), .Q(\values[92] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[91]_reg  (.CK(clk), .E(n_91), .SE(1'b0), 
      .GCK(n_121_28));
   DFF_X1 \values_reg[91][15]  (.D(values[15]), .CK(n_121_28), .Q(
      \values[91] [15]), .QN());
   DFF_X1 \values_reg[91][14]  (.D(values[14]), .CK(n_121_28), .Q(
      \values[91] [14]), .QN());
   DFF_X1 \values_reg[91][13]  (.D(values[13]), .CK(n_121_28), .Q(
      \values[91] [13]), .QN());
   DFF_X1 \values_reg[91][12]  (.D(values[12]), .CK(n_121_28), .Q(
      \values[91] [12]), .QN());
   DFF_X1 \values_reg[91][11]  (.D(values[11]), .CK(n_121_28), .Q(
      \values[91] [11]), .QN());
   DFF_X1 \values_reg[91][10]  (.D(values[10]), .CK(n_121_28), .Q(
      \values[91] [10]), .QN());
   DFF_X1 \values_reg[91][9]  (.D(values[9]), .CK(n_121_28), .Q(\values[91] [9]), 
      .QN());
   DFF_X1 \values_reg[91][8]  (.D(values[8]), .CK(n_121_28), .Q(\values[91] [8]), 
      .QN());
   DFF_X1 \values_reg[91][7]  (.D(values[7]), .CK(n_121_28), .Q(\values[91] [7]), 
      .QN());
   DFF_X1 \values_reg[91][6]  (.D(values[6]), .CK(n_121_28), .Q(\values[91] [6]), 
      .QN());
   DFF_X1 \values_reg[91][5]  (.D(values[5]), .CK(n_121_28), .Q(\values[91] [5]), 
      .QN());
   DFF_X1 \values_reg[91][4]  (.D(values[4]), .CK(n_121_28), .Q(\values[91] [4]), 
      .QN());
   DFF_X1 \values_reg[91][3]  (.D(values[3]), .CK(n_121_28), .Q(\values[91] [3]), 
      .QN());
   DFF_X1 \values_reg[91][2]  (.D(values[2]), .CK(n_121_28), .Q(\values[91] [2]), 
      .QN());
   DFF_X1 \values_reg[91][1]  (.D(values[1]), .CK(n_121_28), .Q(\values[91] [1]), 
      .QN());
   DFF_X1 \values_reg[91][0]  (.D(values[0]), .CK(n_121_28), .Q(\values[91] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[90]_reg  (.CK(clk), .E(n_90), .SE(1'b0), 
      .GCK(n_121_29));
   DFF_X1 \values_reg[90][15]  (.D(values[15]), .CK(n_121_29), .Q(
      \values[90] [15]), .QN());
   DFF_X1 \values_reg[90][14]  (.D(values[14]), .CK(n_121_29), .Q(
      \values[90] [14]), .QN());
   DFF_X1 \values_reg[90][13]  (.D(values[13]), .CK(n_121_29), .Q(
      \values[90] [13]), .QN());
   DFF_X1 \values_reg[90][12]  (.D(values[12]), .CK(n_121_29), .Q(
      \values[90] [12]), .QN());
   DFF_X1 \values_reg[90][11]  (.D(values[11]), .CK(n_121_29), .Q(
      \values[90] [11]), .QN());
   DFF_X1 \values_reg[90][10]  (.D(values[10]), .CK(n_121_29), .Q(
      \values[90] [10]), .QN());
   DFF_X1 \values_reg[90][9]  (.D(values[9]), .CK(n_121_29), .Q(\values[90] [9]), 
      .QN());
   DFF_X1 \values_reg[90][8]  (.D(values[8]), .CK(n_121_29), .Q(\values[90] [8]), 
      .QN());
   DFF_X1 \values_reg[90][7]  (.D(values[7]), .CK(n_121_29), .Q(\values[90] [7]), 
      .QN());
   DFF_X1 \values_reg[90][6]  (.D(values[6]), .CK(n_121_29), .Q(\values[90] [6]), 
      .QN());
   DFF_X1 \values_reg[90][5]  (.D(values[5]), .CK(n_121_29), .Q(\values[90] [5]), 
      .QN());
   DFF_X1 \values_reg[90][4]  (.D(values[4]), .CK(n_121_29), .Q(\values[90] [4]), 
      .QN());
   DFF_X1 \values_reg[90][3]  (.D(values[3]), .CK(n_121_29), .Q(\values[90] [3]), 
      .QN());
   DFF_X1 \values_reg[90][2]  (.D(values[2]), .CK(n_121_29), .Q(\values[90] [2]), 
      .QN());
   DFF_X1 \values_reg[90][1]  (.D(values[1]), .CK(n_121_29), .Q(\values[90] [1]), 
      .QN());
   DFF_X1 \values_reg[90][0]  (.D(values[0]), .CK(n_121_29), .Q(\values[90] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[89]_reg  (.CK(clk), .E(n_89), .SE(1'b0), 
      .GCK(n_121_30));
   DFF_X1 \values_reg[89][15]  (.D(values[15]), .CK(n_121_30), .Q(
      \values[89] [15]), .QN());
   DFF_X1 \values_reg[89][14]  (.D(values[14]), .CK(n_121_30), .Q(
      \values[89] [14]), .QN());
   DFF_X1 \values_reg[89][13]  (.D(values[13]), .CK(n_121_30), .Q(
      \values[89] [13]), .QN());
   DFF_X1 \values_reg[89][12]  (.D(values[12]), .CK(n_121_30), .Q(
      \values[89] [12]), .QN());
   DFF_X1 \values_reg[89][11]  (.D(values[11]), .CK(n_121_30), .Q(
      \values[89] [11]), .QN());
   DFF_X1 \values_reg[89][10]  (.D(values[10]), .CK(n_121_30), .Q(
      \values[89] [10]), .QN());
   DFF_X1 \values_reg[89][9]  (.D(values[9]), .CK(n_121_30), .Q(\values[89] [9]), 
      .QN());
   DFF_X1 \values_reg[89][8]  (.D(values[8]), .CK(n_121_30), .Q(\values[89] [8]), 
      .QN());
   DFF_X1 \values_reg[89][7]  (.D(values[7]), .CK(n_121_30), .Q(\values[89] [7]), 
      .QN());
   DFF_X1 \values_reg[89][6]  (.D(values[6]), .CK(n_121_30), .Q(\values[89] [6]), 
      .QN());
   DFF_X1 \values_reg[89][5]  (.D(values[5]), .CK(n_121_30), .Q(\values[89] [5]), 
      .QN());
   DFF_X1 \values_reg[89][4]  (.D(values[4]), .CK(n_121_30), .Q(\values[89] [4]), 
      .QN());
   DFF_X1 \values_reg[89][3]  (.D(values[3]), .CK(n_121_30), .Q(\values[89] [3]), 
      .QN());
   DFF_X1 \values_reg[89][2]  (.D(values[2]), .CK(n_121_30), .Q(\values[89] [2]), 
      .QN());
   DFF_X1 \values_reg[89][1]  (.D(values[1]), .CK(n_121_30), .Q(\values[89] [1]), 
      .QN());
   DFF_X1 \values_reg[89][0]  (.D(values[0]), .CK(n_121_30), .Q(\values[89] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[88]_reg  (.CK(clk), .E(n_88), .SE(1'b0), 
      .GCK(n_121_31));
   DFF_X1 \values_reg[88][15]  (.D(values[15]), .CK(n_121_31), .Q(
      \values[88] [15]), .QN());
   DFF_X1 \values_reg[88][14]  (.D(values[14]), .CK(n_121_31), .Q(
      \values[88] [14]), .QN());
   DFF_X1 \values_reg[88][13]  (.D(values[13]), .CK(n_121_31), .Q(
      \values[88] [13]), .QN());
   DFF_X1 \values_reg[88][12]  (.D(values[12]), .CK(n_121_31), .Q(
      \values[88] [12]), .QN());
   DFF_X1 \values_reg[88][11]  (.D(values[11]), .CK(n_121_31), .Q(
      \values[88] [11]), .QN());
   DFF_X1 \values_reg[88][10]  (.D(values[10]), .CK(n_121_31), .Q(
      \values[88] [10]), .QN());
   DFF_X1 \values_reg[88][9]  (.D(values[9]), .CK(n_121_31), .Q(\values[88] [9]), 
      .QN());
   DFF_X1 \values_reg[88][8]  (.D(values[8]), .CK(n_121_31), .Q(\values[88] [8]), 
      .QN());
   DFF_X1 \values_reg[88][7]  (.D(values[7]), .CK(n_121_31), .Q(\values[88] [7]), 
      .QN());
   DFF_X1 \values_reg[88][6]  (.D(values[6]), .CK(n_121_31), .Q(\values[88] [6]), 
      .QN());
   DFF_X1 \values_reg[88][5]  (.D(values[5]), .CK(n_121_31), .Q(\values[88] [5]), 
      .QN());
   DFF_X1 \values_reg[88][4]  (.D(values[4]), .CK(n_121_31), .Q(\values[88] [4]), 
      .QN());
   DFF_X1 \values_reg[88][3]  (.D(values[3]), .CK(n_121_31), .Q(\values[88] [3]), 
      .QN());
   DFF_X1 \values_reg[88][2]  (.D(values[2]), .CK(n_121_31), .Q(\values[88] [2]), 
      .QN());
   DFF_X1 \values_reg[88][1]  (.D(values[1]), .CK(n_121_31), .Q(\values[88] [1]), 
      .QN());
   DFF_X1 \values_reg[88][0]  (.D(values[0]), .CK(n_121_31), .Q(\values[88] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[87]_reg  (.CK(clk), .E(n_87), .SE(1'b0), 
      .GCK(n_121_32));
   DFF_X1 \values_reg[87][15]  (.D(values[15]), .CK(n_121_32), .Q(
      \values[87] [15]), .QN());
   DFF_X1 \values_reg[87][14]  (.D(values[14]), .CK(n_121_32), .Q(
      \values[87] [14]), .QN());
   DFF_X1 \values_reg[87][13]  (.D(values[13]), .CK(n_121_32), .Q(
      \values[87] [13]), .QN());
   DFF_X1 \values_reg[87][12]  (.D(values[12]), .CK(n_121_32), .Q(
      \values[87] [12]), .QN());
   DFF_X1 \values_reg[87][11]  (.D(values[11]), .CK(n_121_32), .Q(
      \values[87] [11]), .QN());
   DFF_X1 \values_reg[87][10]  (.D(values[10]), .CK(n_121_32), .Q(
      \values[87] [10]), .QN());
   DFF_X1 \values_reg[87][9]  (.D(values[9]), .CK(n_121_32), .Q(\values[87] [9]), 
      .QN());
   DFF_X1 \values_reg[87][8]  (.D(values[8]), .CK(n_121_32), .Q(\values[87] [8]), 
      .QN());
   DFF_X1 \values_reg[87][7]  (.D(values[7]), .CK(n_121_32), .Q(\values[87] [7]), 
      .QN());
   DFF_X1 \values_reg[87][6]  (.D(values[6]), .CK(n_121_32), .Q(\values[87] [6]), 
      .QN());
   DFF_X1 \values_reg[87][5]  (.D(values[5]), .CK(n_121_32), .Q(\values[87] [5]), 
      .QN());
   DFF_X1 \values_reg[87][4]  (.D(values[4]), .CK(n_121_32), .Q(\values[87] [4]), 
      .QN());
   DFF_X1 \values_reg[87][3]  (.D(values[3]), .CK(n_121_32), .Q(\values[87] [3]), 
      .QN());
   DFF_X1 \values_reg[87][2]  (.D(values[2]), .CK(n_121_32), .Q(\values[87] [2]), 
      .QN());
   DFF_X1 \values_reg[87][1]  (.D(values[1]), .CK(n_121_32), .Q(\values[87] [1]), 
      .QN());
   DFF_X1 \values_reg[87][0]  (.D(values[0]), .CK(n_121_32), .Q(\values[87] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[86]_reg  (.CK(clk), .E(n_86), .SE(1'b0), 
      .GCK(n_121_33));
   DFF_X1 \values_reg[86][15]  (.D(values[15]), .CK(n_121_33), .Q(
      \values[86] [15]), .QN());
   DFF_X1 \values_reg[86][14]  (.D(values[14]), .CK(n_121_33), .Q(
      \values[86] [14]), .QN());
   DFF_X1 \values_reg[86][13]  (.D(values[13]), .CK(n_121_33), .Q(
      \values[86] [13]), .QN());
   DFF_X1 \values_reg[86][12]  (.D(values[12]), .CK(n_121_33), .Q(
      \values[86] [12]), .QN());
   DFF_X1 \values_reg[86][11]  (.D(values[11]), .CK(n_121_33), .Q(
      \values[86] [11]), .QN());
   DFF_X1 \values_reg[86][10]  (.D(values[10]), .CK(n_121_33), .Q(
      \values[86] [10]), .QN());
   DFF_X1 \values_reg[86][9]  (.D(values[9]), .CK(n_121_33), .Q(\values[86] [9]), 
      .QN());
   DFF_X1 \values_reg[86][8]  (.D(values[8]), .CK(n_121_33), .Q(\values[86] [8]), 
      .QN());
   DFF_X1 \values_reg[86][7]  (.D(values[7]), .CK(n_121_33), .Q(\values[86] [7]), 
      .QN());
   DFF_X1 \values_reg[86][6]  (.D(values[6]), .CK(n_121_33), .Q(\values[86] [6]), 
      .QN());
   DFF_X1 \values_reg[86][5]  (.D(values[5]), .CK(n_121_33), .Q(\values[86] [5]), 
      .QN());
   DFF_X1 \values_reg[86][4]  (.D(values[4]), .CK(n_121_33), .Q(\values[86] [4]), 
      .QN());
   DFF_X1 \values_reg[86][3]  (.D(values[3]), .CK(n_121_33), .Q(\values[86] [3]), 
      .QN());
   DFF_X1 \values_reg[86][2]  (.D(values[2]), .CK(n_121_33), .Q(\values[86] [2]), 
      .QN());
   DFF_X1 \values_reg[86][1]  (.D(values[1]), .CK(n_121_33), .Q(\values[86] [1]), 
      .QN());
   DFF_X1 \values_reg[86][0]  (.D(values[0]), .CK(n_121_33), .Q(\values[86] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[85]_reg  (.CK(clk), .E(n_85), .SE(1'b0), 
      .GCK(n_121_34));
   DFF_X1 \values_reg[85][15]  (.D(values[15]), .CK(n_121_34), .Q(
      \values[85] [15]), .QN());
   DFF_X1 \values_reg[85][14]  (.D(values[14]), .CK(n_121_34), .Q(
      \values[85] [14]), .QN());
   DFF_X1 \values_reg[85][13]  (.D(values[13]), .CK(n_121_34), .Q(
      \values[85] [13]), .QN());
   DFF_X1 \values_reg[85][12]  (.D(values[12]), .CK(n_121_34), .Q(
      \values[85] [12]), .QN());
   DFF_X1 \values_reg[85][11]  (.D(values[11]), .CK(n_121_34), .Q(
      \values[85] [11]), .QN());
   DFF_X1 \values_reg[85][10]  (.D(values[10]), .CK(n_121_34), .Q(
      \values[85] [10]), .QN());
   DFF_X1 \values_reg[85][9]  (.D(values[9]), .CK(n_121_34), .Q(\values[85] [9]), 
      .QN());
   DFF_X1 \values_reg[85][8]  (.D(values[8]), .CK(n_121_34), .Q(\values[85] [8]), 
      .QN());
   DFF_X1 \values_reg[85][7]  (.D(values[7]), .CK(n_121_34), .Q(\values[85] [7]), 
      .QN());
   DFF_X1 \values_reg[85][6]  (.D(values[6]), .CK(n_121_34), .Q(\values[85] [6]), 
      .QN());
   DFF_X1 \values_reg[85][5]  (.D(values[5]), .CK(n_121_34), .Q(\values[85] [5]), 
      .QN());
   DFF_X1 \values_reg[85][4]  (.D(values[4]), .CK(n_121_34), .Q(\values[85] [4]), 
      .QN());
   DFF_X1 \values_reg[85][3]  (.D(values[3]), .CK(n_121_34), .Q(\values[85] [3]), 
      .QN());
   DFF_X1 \values_reg[85][2]  (.D(values[2]), .CK(n_121_34), .Q(\values[85] [2]), 
      .QN());
   DFF_X1 \values_reg[85][1]  (.D(values[1]), .CK(n_121_34), .Q(\values[85] [1]), 
      .QN());
   DFF_X1 \values_reg[85][0]  (.D(values[0]), .CK(n_121_34), .Q(\values[85] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[84]_reg  (.CK(clk), .E(n_84), .SE(1'b0), 
      .GCK(n_121_35));
   DFF_X1 \values_reg[84][15]  (.D(values[15]), .CK(n_121_35), .Q(
      \values[84] [15]), .QN());
   DFF_X1 \values_reg[84][14]  (.D(values[14]), .CK(n_121_35), .Q(
      \values[84] [14]), .QN());
   DFF_X1 \values_reg[84][13]  (.D(values[13]), .CK(n_121_35), .Q(
      \values[84] [13]), .QN());
   DFF_X1 \values_reg[84][12]  (.D(values[12]), .CK(n_121_35), .Q(
      \values[84] [12]), .QN());
   DFF_X1 \values_reg[84][11]  (.D(values[11]), .CK(n_121_35), .Q(
      \values[84] [11]), .QN());
   DFF_X1 \values_reg[84][10]  (.D(values[10]), .CK(n_121_35), .Q(
      \values[84] [10]), .QN());
   DFF_X1 \values_reg[84][9]  (.D(values[9]), .CK(n_121_35), .Q(\values[84] [9]), 
      .QN());
   DFF_X1 \values_reg[84][8]  (.D(values[8]), .CK(n_121_35), .Q(\values[84] [8]), 
      .QN());
   DFF_X1 \values_reg[84][7]  (.D(values[7]), .CK(n_121_35), .Q(\values[84] [7]), 
      .QN());
   DFF_X1 \values_reg[84][6]  (.D(values[6]), .CK(n_121_35), .Q(\values[84] [6]), 
      .QN());
   DFF_X1 \values_reg[84][5]  (.D(values[5]), .CK(n_121_35), .Q(\values[84] [5]), 
      .QN());
   DFF_X1 \values_reg[84][4]  (.D(values[4]), .CK(n_121_35), .Q(\values[84] [4]), 
      .QN());
   DFF_X1 \values_reg[84][3]  (.D(values[3]), .CK(n_121_35), .Q(\values[84] [3]), 
      .QN());
   DFF_X1 \values_reg[84][2]  (.D(values[2]), .CK(n_121_35), .Q(\values[84] [2]), 
      .QN());
   DFF_X1 \values_reg[84][1]  (.D(values[1]), .CK(n_121_35), .Q(\values[84] [1]), 
      .QN());
   DFF_X1 \values_reg[84][0]  (.D(values[0]), .CK(n_121_35), .Q(\values[84] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[83]_reg  (.CK(clk), .E(n_83), .SE(1'b0), 
      .GCK(n_121_36));
   DFF_X1 \values_reg[83][15]  (.D(values[15]), .CK(n_121_36), .Q(
      \values[83] [15]), .QN());
   DFF_X1 \values_reg[83][14]  (.D(values[14]), .CK(n_121_36), .Q(
      \values[83] [14]), .QN());
   DFF_X1 \values_reg[83][13]  (.D(values[13]), .CK(n_121_36), .Q(
      \values[83] [13]), .QN());
   DFF_X1 \values_reg[83][12]  (.D(values[12]), .CK(n_121_36), .Q(
      \values[83] [12]), .QN());
   DFF_X1 \values_reg[83][11]  (.D(values[11]), .CK(n_121_36), .Q(
      \values[83] [11]), .QN());
   DFF_X1 \values_reg[83][10]  (.D(values[10]), .CK(n_121_36), .Q(
      \values[83] [10]), .QN());
   DFF_X1 \values_reg[83][9]  (.D(values[9]), .CK(n_121_36), .Q(\values[83] [9]), 
      .QN());
   DFF_X1 \values_reg[83][8]  (.D(values[8]), .CK(n_121_36), .Q(\values[83] [8]), 
      .QN());
   DFF_X1 \values_reg[83][7]  (.D(values[7]), .CK(n_121_36), .Q(\values[83] [7]), 
      .QN());
   DFF_X1 \values_reg[83][6]  (.D(values[6]), .CK(n_121_36), .Q(\values[83] [6]), 
      .QN());
   DFF_X1 \values_reg[83][5]  (.D(values[5]), .CK(n_121_36), .Q(\values[83] [5]), 
      .QN());
   DFF_X1 \values_reg[83][4]  (.D(values[4]), .CK(n_121_36), .Q(\values[83] [4]), 
      .QN());
   DFF_X1 \values_reg[83][3]  (.D(values[3]), .CK(n_121_36), .Q(\values[83] [3]), 
      .QN());
   DFF_X1 \values_reg[83][2]  (.D(values[2]), .CK(n_121_36), .Q(\values[83] [2]), 
      .QN());
   DFF_X1 \values_reg[83][1]  (.D(values[1]), .CK(n_121_36), .Q(\values[83] [1]), 
      .QN());
   DFF_X1 \values_reg[83][0]  (.D(values[0]), .CK(n_121_36), .Q(\values[83] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[82]_reg  (.CK(clk), .E(n_82), .SE(1'b0), 
      .GCK(n_121_37));
   DFF_X1 \values_reg[82][15]  (.D(values[15]), .CK(n_121_37), .Q(
      \values[82] [15]), .QN());
   DFF_X1 \values_reg[82][14]  (.D(values[14]), .CK(n_121_37), .Q(
      \values[82] [14]), .QN());
   DFF_X1 \values_reg[82][13]  (.D(values[13]), .CK(n_121_37), .Q(
      \values[82] [13]), .QN());
   DFF_X1 \values_reg[82][12]  (.D(values[12]), .CK(n_121_37), .Q(
      \values[82] [12]), .QN());
   DFF_X1 \values_reg[82][11]  (.D(values[11]), .CK(n_121_37), .Q(
      \values[82] [11]), .QN());
   DFF_X1 \values_reg[82][10]  (.D(values[10]), .CK(n_121_37), .Q(
      \values[82] [10]), .QN());
   DFF_X1 \values_reg[82][9]  (.D(values[9]), .CK(n_121_37), .Q(\values[82] [9]), 
      .QN());
   DFF_X1 \values_reg[82][8]  (.D(values[8]), .CK(n_121_37), .Q(\values[82] [8]), 
      .QN());
   DFF_X1 \values_reg[82][7]  (.D(values[7]), .CK(n_121_37), .Q(\values[82] [7]), 
      .QN());
   DFF_X1 \values_reg[82][6]  (.D(values[6]), .CK(n_121_37), .Q(\values[82] [6]), 
      .QN());
   DFF_X1 \values_reg[82][5]  (.D(values[5]), .CK(n_121_37), .Q(\values[82] [5]), 
      .QN());
   DFF_X1 \values_reg[82][4]  (.D(values[4]), .CK(n_121_37), .Q(\values[82] [4]), 
      .QN());
   DFF_X1 \values_reg[82][3]  (.D(values[3]), .CK(n_121_37), .Q(\values[82] [3]), 
      .QN());
   DFF_X1 \values_reg[82][2]  (.D(values[2]), .CK(n_121_37), .Q(\values[82] [2]), 
      .QN());
   DFF_X1 \values_reg[82][1]  (.D(values[1]), .CK(n_121_37), .Q(\values[82] [1]), 
      .QN());
   DFF_X1 \values_reg[82][0]  (.D(values[0]), .CK(n_121_37), .Q(\values[82] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[81]_reg  (.CK(clk), .E(n_81), .SE(1'b0), 
      .GCK(n_121_38));
   DFF_X1 \values_reg[81][15]  (.D(values[15]), .CK(n_121_38), .Q(
      \values[81] [15]), .QN());
   DFF_X1 \values_reg[81][14]  (.D(values[14]), .CK(n_121_38), .Q(
      \values[81] [14]), .QN());
   DFF_X1 \values_reg[81][13]  (.D(values[13]), .CK(n_121_38), .Q(
      \values[81] [13]), .QN());
   DFF_X1 \values_reg[81][12]  (.D(values[12]), .CK(n_121_38), .Q(
      \values[81] [12]), .QN());
   DFF_X1 \values_reg[81][11]  (.D(values[11]), .CK(n_121_38), .Q(
      \values[81] [11]), .QN());
   DFF_X1 \values_reg[81][10]  (.D(values[10]), .CK(n_121_38), .Q(
      \values[81] [10]), .QN());
   DFF_X1 \values_reg[81][9]  (.D(values[9]), .CK(n_121_38), .Q(\values[81] [9]), 
      .QN());
   DFF_X1 \values_reg[81][8]  (.D(values[8]), .CK(n_121_38), .Q(\values[81] [8]), 
      .QN());
   DFF_X1 \values_reg[81][7]  (.D(values[7]), .CK(n_121_38), .Q(\values[81] [7]), 
      .QN());
   DFF_X1 \values_reg[81][6]  (.D(values[6]), .CK(n_121_38), .Q(\values[81] [6]), 
      .QN());
   DFF_X1 \values_reg[81][5]  (.D(values[5]), .CK(n_121_38), .Q(\values[81] [5]), 
      .QN());
   DFF_X1 \values_reg[81][4]  (.D(values[4]), .CK(n_121_38), .Q(\values[81] [4]), 
      .QN());
   DFF_X1 \values_reg[81][3]  (.D(values[3]), .CK(n_121_38), .Q(\values[81] [3]), 
      .QN());
   DFF_X1 \values_reg[81][2]  (.D(values[2]), .CK(n_121_38), .Q(\values[81] [2]), 
      .QN());
   DFF_X1 \values_reg[81][1]  (.D(values[1]), .CK(n_121_38), .Q(\values[81] [1]), 
      .QN());
   DFF_X1 \values_reg[81][0]  (.D(values[0]), .CK(n_121_38), .Q(\values[81] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[80]_reg  (.CK(clk), .E(n_80), .SE(1'b0), 
      .GCK(n_121_39));
   DFF_X1 \values_reg[80][15]  (.D(values[15]), .CK(n_121_39), .Q(
      \values[80] [15]), .QN());
   DFF_X1 \values_reg[80][14]  (.D(values[14]), .CK(n_121_39), .Q(
      \values[80] [14]), .QN());
   DFF_X1 \values_reg[80][13]  (.D(values[13]), .CK(n_121_39), .Q(
      \values[80] [13]), .QN());
   DFF_X1 \values_reg[80][12]  (.D(values[12]), .CK(n_121_39), .Q(
      \values[80] [12]), .QN());
   DFF_X1 \values_reg[80][11]  (.D(values[11]), .CK(n_121_39), .Q(
      \values[80] [11]), .QN());
   DFF_X1 \values_reg[80][10]  (.D(values[10]), .CK(n_121_39), .Q(
      \values[80] [10]), .QN());
   DFF_X1 \values_reg[80][9]  (.D(values[9]), .CK(n_121_39), .Q(\values[80] [9]), 
      .QN());
   DFF_X1 \values_reg[80][8]  (.D(values[8]), .CK(n_121_39), .Q(\values[80] [8]), 
      .QN());
   DFF_X1 \values_reg[80][7]  (.D(values[7]), .CK(n_121_39), .Q(\values[80] [7]), 
      .QN());
   DFF_X1 \values_reg[80][6]  (.D(values[6]), .CK(n_121_39), .Q(\values[80] [6]), 
      .QN());
   DFF_X1 \values_reg[80][5]  (.D(values[5]), .CK(n_121_39), .Q(\values[80] [5]), 
      .QN());
   DFF_X1 \values_reg[80][4]  (.D(values[4]), .CK(n_121_39), .Q(\values[80] [4]), 
      .QN());
   DFF_X1 \values_reg[80][3]  (.D(values[3]), .CK(n_121_39), .Q(\values[80] [3]), 
      .QN());
   DFF_X1 \values_reg[80][2]  (.D(values[2]), .CK(n_121_39), .Q(\values[80] [2]), 
      .QN());
   DFF_X1 \values_reg[80][1]  (.D(values[1]), .CK(n_121_39), .Q(\values[80] [1]), 
      .QN());
   DFF_X1 \values_reg[80][0]  (.D(values[0]), .CK(n_121_39), .Q(\values[80] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[79]_reg  (.CK(clk), .E(n_79), .SE(1'b0), 
      .GCK(n_121_40));
   DFF_X1 \values_reg[79][15]  (.D(values[15]), .CK(n_121_40), .Q(
      \values[79] [15]), .QN());
   DFF_X1 \values_reg[79][14]  (.D(values[14]), .CK(n_121_40), .Q(
      \values[79] [14]), .QN());
   DFF_X1 \values_reg[79][13]  (.D(values[13]), .CK(n_121_40), .Q(
      \values[79] [13]), .QN());
   DFF_X1 \values_reg[79][12]  (.D(values[12]), .CK(n_121_40), .Q(
      \values[79] [12]), .QN());
   DFF_X1 \values_reg[79][11]  (.D(values[11]), .CK(n_121_40), .Q(
      \values[79] [11]), .QN());
   DFF_X1 \values_reg[79][10]  (.D(values[10]), .CK(n_121_40), .Q(
      \values[79] [10]), .QN());
   DFF_X1 \values_reg[79][9]  (.D(values[9]), .CK(n_121_40), .Q(\values[79] [9]), 
      .QN());
   DFF_X1 \values_reg[79][8]  (.D(values[8]), .CK(n_121_40), .Q(\values[79] [8]), 
      .QN());
   DFF_X1 \values_reg[79][7]  (.D(values[7]), .CK(n_121_40), .Q(\values[79] [7]), 
      .QN());
   DFF_X1 \values_reg[79][6]  (.D(values[6]), .CK(n_121_40), .Q(\values[79] [6]), 
      .QN());
   DFF_X1 \values_reg[79][5]  (.D(values[5]), .CK(n_121_40), .Q(\values[79] [5]), 
      .QN());
   DFF_X1 \values_reg[79][4]  (.D(values[4]), .CK(n_121_40), .Q(\values[79] [4]), 
      .QN());
   DFF_X1 \values_reg[79][3]  (.D(values[3]), .CK(n_121_40), .Q(\values[79] [3]), 
      .QN());
   DFF_X1 \values_reg[79][2]  (.D(values[2]), .CK(n_121_40), .Q(\values[79] [2]), 
      .QN());
   DFF_X1 \values_reg[79][1]  (.D(values[1]), .CK(n_121_40), .Q(\values[79] [1]), 
      .QN());
   DFF_X1 \values_reg[79][0]  (.D(values[0]), .CK(n_121_40), .Q(\values[79] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[78]_reg  (.CK(clk), .E(n_78), .SE(1'b0), 
      .GCK(n_121_41));
   DFF_X1 \values_reg[78][15]  (.D(values[15]), .CK(n_121_41), .Q(
      \values[78] [15]), .QN());
   DFF_X1 \values_reg[78][14]  (.D(values[14]), .CK(n_121_41), .Q(
      \values[78] [14]), .QN());
   DFF_X1 \values_reg[78][13]  (.D(values[13]), .CK(n_121_41), .Q(
      \values[78] [13]), .QN());
   DFF_X1 \values_reg[78][12]  (.D(values[12]), .CK(n_121_41), .Q(
      \values[78] [12]), .QN());
   DFF_X1 \values_reg[78][11]  (.D(values[11]), .CK(n_121_41), .Q(
      \values[78] [11]), .QN());
   DFF_X1 \values_reg[78][10]  (.D(values[10]), .CK(n_121_41), .Q(
      \values[78] [10]), .QN());
   DFF_X1 \values_reg[78][9]  (.D(values[9]), .CK(n_121_41), .Q(\values[78] [9]), 
      .QN());
   DFF_X1 \values_reg[78][8]  (.D(values[8]), .CK(n_121_41), .Q(\values[78] [8]), 
      .QN());
   DFF_X1 \values_reg[78][7]  (.D(values[7]), .CK(n_121_41), .Q(\values[78] [7]), 
      .QN());
   DFF_X1 \values_reg[78][6]  (.D(values[6]), .CK(n_121_41), .Q(\values[78] [6]), 
      .QN());
   DFF_X1 \values_reg[78][5]  (.D(values[5]), .CK(n_121_41), .Q(\values[78] [5]), 
      .QN());
   DFF_X1 \values_reg[78][4]  (.D(values[4]), .CK(n_121_41), .Q(\values[78] [4]), 
      .QN());
   DFF_X1 \values_reg[78][3]  (.D(values[3]), .CK(n_121_41), .Q(\values[78] [3]), 
      .QN());
   DFF_X1 \values_reg[78][2]  (.D(values[2]), .CK(n_121_41), .Q(\values[78] [2]), 
      .QN());
   DFF_X1 \values_reg[78][1]  (.D(values[1]), .CK(n_121_41), .Q(\values[78] [1]), 
      .QN());
   DFF_X1 \values_reg[78][0]  (.D(values[0]), .CK(n_121_41), .Q(\values[78] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[77]_reg  (.CK(clk), .E(n_77), .SE(1'b0), 
      .GCK(n_121_42));
   DFF_X1 \values_reg[77][15]  (.D(values[15]), .CK(n_121_42), .Q(
      \values[77] [15]), .QN());
   DFF_X1 \values_reg[77][14]  (.D(values[14]), .CK(n_121_42), .Q(
      \values[77] [14]), .QN());
   DFF_X1 \values_reg[77][13]  (.D(values[13]), .CK(n_121_42), .Q(
      \values[77] [13]), .QN());
   DFF_X1 \values_reg[77][12]  (.D(values[12]), .CK(n_121_42), .Q(
      \values[77] [12]), .QN());
   DFF_X1 \values_reg[77][11]  (.D(values[11]), .CK(n_121_42), .Q(
      \values[77] [11]), .QN());
   DFF_X1 \values_reg[77][10]  (.D(values[10]), .CK(n_121_42), .Q(
      \values[77] [10]), .QN());
   DFF_X1 \values_reg[77][9]  (.D(values[9]), .CK(n_121_42), .Q(\values[77] [9]), 
      .QN());
   DFF_X1 \values_reg[77][8]  (.D(values[8]), .CK(n_121_42), .Q(\values[77] [8]), 
      .QN());
   DFF_X1 \values_reg[77][7]  (.D(values[7]), .CK(n_121_42), .Q(\values[77] [7]), 
      .QN());
   DFF_X1 \values_reg[77][6]  (.D(values[6]), .CK(n_121_42), .Q(\values[77] [6]), 
      .QN());
   DFF_X1 \values_reg[77][5]  (.D(values[5]), .CK(n_121_42), .Q(\values[77] [5]), 
      .QN());
   DFF_X1 \values_reg[77][4]  (.D(values[4]), .CK(n_121_42), .Q(\values[77] [4]), 
      .QN());
   DFF_X1 \values_reg[77][3]  (.D(values[3]), .CK(n_121_42), .Q(\values[77] [3]), 
      .QN());
   DFF_X1 \values_reg[77][2]  (.D(values[2]), .CK(n_121_42), .Q(\values[77] [2]), 
      .QN());
   DFF_X1 \values_reg[77][1]  (.D(values[1]), .CK(n_121_42), .Q(\values[77] [1]), 
      .QN());
   DFF_X1 \values_reg[77][0]  (.D(values[0]), .CK(n_121_42), .Q(\values[77] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[76]_reg  (.CK(clk), .E(n_76), .SE(1'b0), 
      .GCK(n_121_43));
   DFF_X1 \values_reg[76][15]  (.D(values[15]), .CK(n_121_43), .Q(
      \values[76] [15]), .QN());
   DFF_X1 \values_reg[76][14]  (.D(values[14]), .CK(n_121_43), .Q(
      \values[76] [14]), .QN());
   DFF_X1 \values_reg[76][13]  (.D(values[13]), .CK(n_121_43), .Q(
      \values[76] [13]), .QN());
   DFF_X1 \values_reg[76][12]  (.D(values[12]), .CK(n_121_43), .Q(
      \values[76] [12]), .QN());
   DFF_X1 \values_reg[76][11]  (.D(values[11]), .CK(n_121_43), .Q(
      \values[76] [11]), .QN());
   DFF_X1 \values_reg[76][10]  (.D(values[10]), .CK(n_121_43), .Q(
      \values[76] [10]), .QN());
   DFF_X1 \values_reg[76][9]  (.D(values[9]), .CK(n_121_43), .Q(\values[76] [9]), 
      .QN());
   DFF_X1 \values_reg[76][8]  (.D(values[8]), .CK(n_121_43), .Q(\values[76] [8]), 
      .QN());
   DFF_X1 \values_reg[76][7]  (.D(values[7]), .CK(n_121_43), .Q(\values[76] [7]), 
      .QN());
   DFF_X1 \values_reg[76][6]  (.D(values[6]), .CK(n_121_43), .Q(\values[76] [6]), 
      .QN());
   DFF_X1 \values_reg[76][5]  (.D(values[5]), .CK(n_121_43), .Q(\values[76] [5]), 
      .QN());
   DFF_X1 \values_reg[76][4]  (.D(values[4]), .CK(n_121_43), .Q(\values[76] [4]), 
      .QN());
   DFF_X1 \values_reg[76][3]  (.D(values[3]), .CK(n_121_43), .Q(\values[76] [3]), 
      .QN());
   DFF_X1 \values_reg[76][2]  (.D(values[2]), .CK(n_121_43), .Q(\values[76] [2]), 
      .QN());
   DFF_X1 \values_reg[76][1]  (.D(values[1]), .CK(n_121_43), .Q(\values[76] [1]), 
      .QN());
   DFF_X1 \values_reg[76][0]  (.D(values[0]), .CK(n_121_43), .Q(\values[76] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[75]_reg  (.CK(clk), .E(n_75), .SE(1'b0), 
      .GCK(n_121_44));
   DFF_X1 \values_reg[75][15]  (.D(values[15]), .CK(n_121_44), .Q(
      \values[75] [15]), .QN());
   DFF_X1 \values_reg[75][14]  (.D(values[14]), .CK(n_121_44), .Q(
      \values[75] [14]), .QN());
   DFF_X1 \values_reg[75][13]  (.D(values[13]), .CK(n_121_44), .Q(
      \values[75] [13]), .QN());
   DFF_X1 \values_reg[75][12]  (.D(values[12]), .CK(n_121_44), .Q(
      \values[75] [12]), .QN());
   DFF_X1 \values_reg[75][11]  (.D(values[11]), .CK(n_121_44), .Q(
      \values[75] [11]), .QN());
   DFF_X1 \values_reg[75][10]  (.D(values[10]), .CK(n_121_44), .Q(
      \values[75] [10]), .QN());
   DFF_X1 \values_reg[75][9]  (.D(values[9]), .CK(n_121_44), .Q(\values[75] [9]), 
      .QN());
   DFF_X1 \values_reg[75][8]  (.D(values[8]), .CK(n_121_44), .Q(\values[75] [8]), 
      .QN());
   DFF_X1 \values_reg[75][7]  (.D(values[7]), .CK(n_121_44), .Q(\values[75] [7]), 
      .QN());
   DFF_X1 \values_reg[75][6]  (.D(values[6]), .CK(n_121_44), .Q(\values[75] [6]), 
      .QN());
   DFF_X1 \values_reg[75][5]  (.D(values[5]), .CK(n_121_44), .Q(\values[75] [5]), 
      .QN());
   DFF_X1 \values_reg[75][4]  (.D(values[4]), .CK(n_121_44), .Q(\values[75] [4]), 
      .QN());
   DFF_X1 \values_reg[75][3]  (.D(values[3]), .CK(n_121_44), .Q(\values[75] [3]), 
      .QN());
   DFF_X1 \values_reg[75][2]  (.D(values[2]), .CK(n_121_44), .Q(\values[75] [2]), 
      .QN());
   DFF_X1 \values_reg[75][1]  (.D(values[1]), .CK(n_121_44), .Q(\values[75] [1]), 
      .QN());
   DFF_X1 \values_reg[75][0]  (.D(values[0]), .CK(n_121_44), .Q(\values[75] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[74]_reg  (.CK(clk), .E(n_74), .SE(1'b0), 
      .GCK(n_121_45));
   DFF_X1 \values_reg[74][15]  (.D(values[15]), .CK(n_121_45), .Q(
      \values[74] [15]), .QN());
   DFF_X1 \values_reg[74][14]  (.D(values[14]), .CK(n_121_45), .Q(
      \values[74] [14]), .QN());
   DFF_X1 \values_reg[74][13]  (.D(values[13]), .CK(n_121_45), .Q(
      \values[74] [13]), .QN());
   DFF_X1 \values_reg[74][12]  (.D(values[12]), .CK(n_121_45), .Q(
      \values[74] [12]), .QN());
   DFF_X1 \values_reg[74][11]  (.D(values[11]), .CK(n_121_45), .Q(
      \values[74] [11]), .QN());
   DFF_X1 \values_reg[74][10]  (.D(values[10]), .CK(n_121_45), .Q(
      \values[74] [10]), .QN());
   DFF_X1 \values_reg[74][9]  (.D(values[9]), .CK(n_121_45), .Q(\values[74] [9]), 
      .QN());
   DFF_X1 \values_reg[74][8]  (.D(values[8]), .CK(n_121_45), .Q(\values[74] [8]), 
      .QN());
   DFF_X1 \values_reg[74][7]  (.D(values[7]), .CK(n_121_45), .Q(\values[74] [7]), 
      .QN());
   DFF_X1 \values_reg[74][6]  (.D(values[6]), .CK(n_121_45), .Q(\values[74] [6]), 
      .QN());
   DFF_X1 \values_reg[74][5]  (.D(values[5]), .CK(n_121_45), .Q(\values[74] [5]), 
      .QN());
   DFF_X1 \values_reg[74][4]  (.D(values[4]), .CK(n_121_45), .Q(\values[74] [4]), 
      .QN());
   DFF_X1 \values_reg[74][3]  (.D(values[3]), .CK(n_121_45), .Q(\values[74] [3]), 
      .QN());
   DFF_X1 \values_reg[74][2]  (.D(values[2]), .CK(n_121_45), .Q(\values[74] [2]), 
      .QN());
   DFF_X1 \values_reg[74][1]  (.D(values[1]), .CK(n_121_45), .Q(\values[74] [1]), 
      .QN());
   DFF_X1 \values_reg[74][0]  (.D(values[0]), .CK(n_121_45), .Q(\values[74] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[73]_reg  (.CK(clk), .E(n_73), .SE(1'b0), 
      .GCK(n_121_46));
   DFF_X1 \values_reg[73][15]  (.D(values[15]), .CK(n_121_46), .Q(
      \values[73] [15]), .QN());
   DFF_X1 \values_reg[73][14]  (.D(values[14]), .CK(n_121_46), .Q(
      \values[73] [14]), .QN());
   DFF_X1 \values_reg[73][13]  (.D(values[13]), .CK(n_121_46), .Q(
      \values[73] [13]), .QN());
   DFF_X1 \values_reg[73][12]  (.D(values[12]), .CK(n_121_46), .Q(
      \values[73] [12]), .QN());
   DFF_X1 \values_reg[73][11]  (.D(values[11]), .CK(n_121_46), .Q(
      \values[73] [11]), .QN());
   DFF_X1 \values_reg[73][10]  (.D(values[10]), .CK(n_121_46), .Q(
      \values[73] [10]), .QN());
   DFF_X1 \values_reg[73][9]  (.D(values[9]), .CK(n_121_46), .Q(\values[73] [9]), 
      .QN());
   DFF_X1 \values_reg[73][8]  (.D(values[8]), .CK(n_121_46), .Q(\values[73] [8]), 
      .QN());
   DFF_X1 \values_reg[73][7]  (.D(values[7]), .CK(n_121_46), .Q(\values[73] [7]), 
      .QN());
   DFF_X1 \values_reg[73][6]  (.D(values[6]), .CK(n_121_46), .Q(\values[73] [6]), 
      .QN());
   DFF_X1 \values_reg[73][5]  (.D(values[5]), .CK(n_121_46), .Q(\values[73] [5]), 
      .QN());
   DFF_X1 \values_reg[73][4]  (.D(values[4]), .CK(n_121_46), .Q(\values[73] [4]), 
      .QN());
   DFF_X1 \values_reg[73][3]  (.D(values[3]), .CK(n_121_46), .Q(\values[73] [3]), 
      .QN());
   DFF_X1 \values_reg[73][2]  (.D(values[2]), .CK(n_121_46), .Q(\values[73] [2]), 
      .QN());
   DFF_X1 \values_reg[73][1]  (.D(values[1]), .CK(n_121_46), .Q(\values[73] [1]), 
      .QN());
   DFF_X1 \values_reg[73][0]  (.D(values[0]), .CK(n_121_46), .Q(\values[73] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[72]_reg  (.CK(clk), .E(n_72), .SE(1'b0), 
      .GCK(n_121_47));
   DFF_X1 \values_reg[72][15]  (.D(values[15]), .CK(n_121_47), .Q(
      \values[72] [15]), .QN());
   DFF_X1 \values_reg[72][14]  (.D(values[14]), .CK(n_121_47), .Q(
      \values[72] [14]), .QN());
   DFF_X1 \values_reg[72][13]  (.D(values[13]), .CK(n_121_47), .Q(
      \values[72] [13]), .QN());
   DFF_X1 \values_reg[72][12]  (.D(values[12]), .CK(n_121_47), .Q(
      \values[72] [12]), .QN());
   DFF_X1 \values_reg[72][11]  (.D(values[11]), .CK(n_121_47), .Q(
      \values[72] [11]), .QN());
   DFF_X1 \values_reg[72][10]  (.D(values[10]), .CK(n_121_47), .Q(
      \values[72] [10]), .QN());
   DFF_X1 \values_reg[72][9]  (.D(values[9]), .CK(n_121_47), .Q(\values[72] [9]), 
      .QN());
   DFF_X1 \values_reg[72][8]  (.D(values[8]), .CK(n_121_47), .Q(\values[72] [8]), 
      .QN());
   DFF_X1 \values_reg[72][7]  (.D(values[7]), .CK(n_121_47), .Q(\values[72] [7]), 
      .QN());
   DFF_X1 \values_reg[72][6]  (.D(values[6]), .CK(n_121_47), .Q(\values[72] [6]), 
      .QN());
   DFF_X1 \values_reg[72][5]  (.D(values[5]), .CK(n_121_47), .Q(\values[72] [5]), 
      .QN());
   DFF_X1 \values_reg[72][4]  (.D(values[4]), .CK(n_121_47), .Q(\values[72] [4]), 
      .QN());
   DFF_X1 \values_reg[72][3]  (.D(values[3]), .CK(n_121_47), .Q(\values[72] [3]), 
      .QN());
   DFF_X1 \values_reg[72][2]  (.D(values[2]), .CK(n_121_47), .Q(\values[72] [2]), 
      .QN());
   DFF_X1 \values_reg[72][1]  (.D(values[1]), .CK(n_121_47), .Q(\values[72] [1]), 
      .QN());
   DFF_X1 \values_reg[72][0]  (.D(values[0]), .CK(n_121_47), .Q(\values[72] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[71]_reg  (.CK(clk), .E(n_71), .SE(1'b0), 
      .GCK(n_121_48));
   DFF_X1 \values_reg[71][15]  (.D(values[15]), .CK(n_121_48), .Q(
      \values[71] [15]), .QN());
   DFF_X1 \values_reg[71][14]  (.D(values[14]), .CK(n_121_48), .Q(
      \values[71] [14]), .QN());
   DFF_X1 \values_reg[71][13]  (.D(values[13]), .CK(n_121_48), .Q(
      \values[71] [13]), .QN());
   DFF_X1 \values_reg[71][12]  (.D(values[12]), .CK(n_121_48), .Q(
      \values[71] [12]), .QN());
   DFF_X1 \values_reg[71][11]  (.D(values[11]), .CK(n_121_48), .Q(
      \values[71] [11]), .QN());
   DFF_X1 \values_reg[71][10]  (.D(values[10]), .CK(n_121_48), .Q(
      \values[71] [10]), .QN());
   DFF_X1 \values_reg[71][9]  (.D(values[9]), .CK(n_121_48), .Q(\values[71] [9]), 
      .QN());
   DFF_X1 \values_reg[71][8]  (.D(values[8]), .CK(n_121_48), .Q(\values[71] [8]), 
      .QN());
   DFF_X1 \values_reg[71][7]  (.D(values[7]), .CK(n_121_48), .Q(\values[71] [7]), 
      .QN());
   DFF_X1 \values_reg[71][6]  (.D(values[6]), .CK(n_121_48), .Q(\values[71] [6]), 
      .QN());
   DFF_X1 \values_reg[71][5]  (.D(values[5]), .CK(n_121_48), .Q(\values[71] [5]), 
      .QN());
   DFF_X1 \values_reg[71][4]  (.D(values[4]), .CK(n_121_48), .Q(\values[71] [4]), 
      .QN());
   DFF_X1 \values_reg[71][3]  (.D(values[3]), .CK(n_121_48), .Q(\values[71] [3]), 
      .QN());
   DFF_X1 \values_reg[71][2]  (.D(values[2]), .CK(n_121_48), .Q(\values[71] [2]), 
      .QN());
   DFF_X1 \values_reg[71][1]  (.D(values[1]), .CK(n_121_48), .Q(\values[71] [1]), 
      .QN());
   DFF_X1 \values_reg[71][0]  (.D(values[0]), .CK(n_121_48), .Q(\values[71] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[70]_reg  (.CK(clk), .E(n_70), .SE(1'b0), 
      .GCK(n_121_49));
   DFF_X1 \values_reg[70][15]  (.D(values[15]), .CK(n_121_49), .Q(
      \values[70] [15]), .QN());
   DFF_X1 \values_reg[70][14]  (.D(values[14]), .CK(n_121_49), .Q(
      \values[70] [14]), .QN());
   DFF_X1 \values_reg[70][13]  (.D(values[13]), .CK(n_121_49), .Q(
      \values[70] [13]), .QN());
   DFF_X1 \values_reg[70][12]  (.D(values[12]), .CK(n_121_49), .Q(
      \values[70] [12]), .QN());
   DFF_X1 \values_reg[70][11]  (.D(values[11]), .CK(n_121_49), .Q(
      \values[70] [11]), .QN());
   DFF_X1 \values_reg[70][10]  (.D(values[10]), .CK(n_121_49), .Q(
      \values[70] [10]), .QN());
   DFF_X1 \values_reg[70][9]  (.D(values[9]), .CK(n_121_49), .Q(\values[70] [9]), 
      .QN());
   DFF_X1 \values_reg[70][8]  (.D(values[8]), .CK(n_121_49), .Q(\values[70] [8]), 
      .QN());
   DFF_X1 \values_reg[70][7]  (.D(values[7]), .CK(n_121_49), .Q(\values[70] [7]), 
      .QN());
   DFF_X1 \values_reg[70][6]  (.D(values[6]), .CK(n_121_49), .Q(\values[70] [6]), 
      .QN());
   DFF_X1 \values_reg[70][5]  (.D(values[5]), .CK(n_121_49), .Q(\values[70] [5]), 
      .QN());
   DFF_X1 \values_reg[70][4]  (.D(values[4]), .CK(n_121_49), .Q(\values[70] [4]), 
      .QN());
   DFF_X1 \values_reg[70][3]  (.D(values[3]), .CK(n_121_49), .Q(\values[70] [3]), 
      .QN());
   DFF_X1 \values_reg[70][2]  (.D(values[2]), .CK(n_121_49), .Q(\values[70] [2]), 
      .QN());
   DFF_X1 \values_reg[70][1]  (.D(values[1]), .CK(n_121_49), .Q(\values[70] [1]), 
      .QN());
   DFF_X1 \values_reg[70][0]  (.D(values[0]), .CK(n_121_49), .Q(\values[70] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[69]_reg  (.CK(clk), .E(n_69), .SE(1'b0), 
      .GCK(n_121_50));
   DFF_X1 \values_reg[69][15]  (.D(values[15]), .CK(n_121_50), .Q(
      \values[69] [15]), .QN());
   DFF_X1 \values_reg[69][14]  (.D(values[14]), .CK(n_121_50), .Q(
      \values[69] [14]), .QN());
   DFF_X1 \values_reg[69][13]  (.D(values[13]), .CK(n_121_50), .Q(
      \values[69] [13]), .QN());
   DFF_X1 \values_reg[69][12]  (.D(values[12]), .CK(n_121_50), .Q(
      \values[69] [12]), .QN());
   DFF_X1 \values_reg[69][11]  (.D(values[11]), .CK(n_121_50), .Q(
      \values[69] [11]), .QN());
   DFF_X1 \values_reg[69][10]  (.D(values[10]), .CK(n_121_50), .Q(
      \values[69] [10]), .QN());
   DFF_X1 \values_reg[69][9]  (.D(values[9]), .CK(n_121_50), .Q(\values[69] [9]), 
      .QN());
   DFF_X1 \values_reg[69][8]  (.D(values[8]), .CK(n_121_50), .Q(\values[69] [8]), 
      .QN());
   DFF_X1 \values_reg[69][7]  (.D(values[7]), .CK(n_121_50), .Q(\values[69] [7]), 
      .QN());
   DFF_X1 \values_reg[69][6]  (.D(values[6]), .CK(n_121_50), .Q(\values[69] [6]), 
      .QN());
   DFF_X1 \values_reg[69][5]  (.D(values[5]), .CK(n_121_50), .Q(\values[69] [5]), 
      .QN());
   DFF_X1 \values_reg[69][4]  (.D(values[4]), .CK(n_121_50), .Q(\values[69] [4]), 
      .QN());
   DFF_X1 \values_reg[69][3]  (.D(values[3]), .CK(n_121_50), .Q(\values[69] [3]), 
      .QN());
   DFF_X1 \values_reg[69][2]  (.D(values[2]), .CK(n_121_50), .Q(\values[69] [2]), 
      .QN());
   DFF_X1 \values_reg[69][1]  (.D(values[1]), .CK(n_121_50), .Q(\values[69] [1]), 
      .QN());
   DFF_X1 \values_reg[69][0]  (.D(values[0]), .CK(n_121_50), .Q(\values[69] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[68]_reg  (.CK(clk), .E(n_68), .SE(1'b0), 
      .GCK(n_121_51));
   DFF_X1 \values_reg[68][15]  (.D(values[15]), .CK(n_121_51), .Q(
      \values[68] [15]), .QN());
   DFF_X1 \values_reg[68][14]  (.D(values[14]), .CK(n_121_51), .Q(
      \values[68] [14]), .QN());
   DFF_X1 \values_reg[68][13]  (.D(values[13]), .CK(n_121_51), .Q(
      \values[68] [13]), .QN());
   DFF_X1 \values_reg[68][12]  (.D(values[12]), .CK(n_121_51), .Q(
      \values[68] [12]), .QN());
   DFF_X1 \values_reg[68][11]  (.D(values[11]), .CK(n_121_51), .Q(
      \values[68] [11]), .QN());
   DFF_X1 \values_reg[68][10]  (.D(values[10]), .CK(n_121_51), .Q(
      \values[68] [10]), .QN());
   DFF_X1 \values_reg[68][9]  (.D(values[9]), .CK(n_121_51), .Q(\values[68] [9]), 
      .QN());
   DFF_X1 \values_reg[68][8]  (.D(values[8]), .CK(n_121_51), .Q(\values[68] [8]), 
      .QN());
   DFF_X1 \values_reg[68][7]  (.D(values[7]), .CK(n_121_51), .Q(\values[68] [7]), 
      .QN());
   DFF_X1 \values_reg[68][6]  (.D(values[6]), .CK(n_121_51), .Q(\values[68] [6]), 
      .QN());
   DFF_X1 \values_reg[68][5]  (.D(values[5]), .CK(n_121_51), .Q(\values[68] [5]), 
      .QN());
   DFF_X1 \values_reg[68][4]  (.D(values[4]), .CK(n_121_51), .Q(\values[68] [4]), 
      .QN());
   DFF_X1 \values_reg[68][3]  (.D(values[3]), .CK(n_121_51), .Q(\values[68] [3]), 
      .QN());
   DFF_X1 \values_reg[68][2]  (.D(values[2]), .CK(n_121_51), .Q(\values[68] [2]), 
      .QN());
   DFF_X1 \values_reg[68][1]  (.D(values[1]), .CK(n_121_51), .Q(\values[68] [1]), 
      .QN());
   DFF_X1 \values_reg[68][0]  (.D(values[0]), .CK(n_121_51), .Q(\values[68] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[67]_reg  (.CK(clk), .E(n_67), .SE(1'b0), 
      .GCK(n_121_52));
   DFF_X1 \values_reg[67][15]  (.D(values[15]), .CK(n_121_52), .Q(
      \values[67] [15]), .QN());
   DFF_X1 \values_reg[67][14]  (.D(values[14]), .CK(n_121_52), .Q(
      \values[67] [14]), .QN());
   DFF_X1 \values_reg[67][13]  (.D(values[13]), .CK(n_121_52), .Q(
      \values[67] [13]), .QN());
   DFF_X1 \values_reg[67][12]  (.D(values[12]), .CK(n_121_52), .Q(
      \values[67] [12]), .QN());
   DFF_X1 \values_reg[67][11]  (.D(values[11]), .CK(n_121_52), .Q(
      \values[67] [11]), .QN());
   DFF_X1 \values_reg[67][10]  (.D(values[10]), .CK(n_121_52), .Q(
      \values[67] [10]), .QN());
   DFF_X1 \values_reg[67][9]  (.D(values[9]), .CK(n_121_52), .Q(\values[67] [9]), 
      .QN());
   DFF_X1 \values_reg[67][8]  (.D(values[8]), .CK(n_121_52), .Q(\values[67] [8]), 
      .QN());
   DFF_X1 \values_reg[67][7]  (.D(values[7]), .CK(n_121_52), .Q(\values[67] [7]), 
      .QN());
   DFF_X1 \values_reg[67][6]  (.D(values[6]), .CK(n_121_52), .Q(\values[67] [6]), 
      .QN());
   DFF_X1 \values_reg[67][5]  (.D(values[5]), .CK(n_121_52), .Q(\values[67] [5]), 
      .QN());
   DFF_X1 \values_reg[67][4]  (.D(values[4]), .CK(n_121_52), .Q(\values[67] [4]), 
      .QN());
   DFF_X1 \values_reg[67][3]  (.D(values[3]), .CK(n_121_52), .Q(\values[67] [3]), 
      .QN());
   DFF_X1 \values_reg[67][2]  (.D(values[2]), .CK(n_121_52), .Q(\values[67] [2]), 
      .QN());
   DFF_X1 \values_reg[67][1]  (.D(values[1]), .CK(n_121_52), .Q(\values[67] [1]), 
      .QN());
   DFF_X1 \values_reg[67][0]  (.D(values[0]), .CK(n_121_52), .Q(\values[67] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[66]_reg  (.CK(clk), .E(n_66), .SE(1'b0), 
      .GCK(n_121_53));
   DFF_X1 \values_reg[66][15]  (.D(values[15]), .CK(n_121_53), .Q(
      \values[66] [15]), .QN());
   DFF_X1 \values_reg[66][14]  (.D(values[14]), .CK(n_121_53), .Q(
      \values[66] [14]), .QN());
   DFF_X1 \values_reg[66][13]  (.D(values[13]), .CK(n_121_53), .Q(
      \values[66] [13]), .QN());
   DFF_X1 \values_reg[66][12]  (.D(values[12]), .CK(n_121_53), .Q(
      \values[66] [12]), .QN());
   DFF_X1 \values_reg[66][11]  (.D(values[11]), .CK(n_121_53), .Q(
      \values[66] [11]), .QN());
   DFF_X1 \values_reg[66][10]  (.D(values[10]), .CK(n_121_53), .Q(
      \values[66] [10]), .QN());
   DFF_X1 \values_reg[66][9]  (.D(values[9]), .CK(n_121_53), .Q(\values[66] [9]), 
      .QN());
   DFF_X1 \values_reg[66][8]  (.D(values[8]), .CK(n_121_53), .Q(\values[66] [8]), 
      .QN());
   DFF_X1 \values_reg[66][7]  (.D(values[7]), .CK(n_121_53), .Q(\values[66] [7]), 
      .QN());
   DFF_X1 \values_reg[66][6]  (.D(values[6]), .CK(n_121_53), .Q(\values[66] [6]), 
      .QN());
   DFF_X1 \values_reg[66][5]  (.D(values[5]), .CK(n_121_53), .Q(\values[66] [5]), 
      .QN());
   DFF_X1 \values_reg[66][4]  (.D(values[4]), .CK(n_121_53), .Q(\values[66] [4]), 
      .QN());
   DFF_X1 \values_reg[66][3]  (.D(values[3]), .CK(n_121_53), .Q(\values[66] [3]), 
      .QN());
   DFF_X1 \values_reg[66][2]  (.D(values[2]), .CK(n_121_53), .Q(\values[66] [2]), 
      .QN());
   DFF_X1 \values_reg[66][1]  (.D(values[1]), .CK(n_121_53), .Q(\values[66] [1]), 
      .QN());
   DFF_X1 \values_reg[66][0]  (.D(values[0]), .CK(n_121_53), .Q(\values[66] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[65]_reg  (.CK(clk), .E(n_65), .SE(1'b0), 
      .GCK(n_121_54));
   DFF_X1 \values_reg[65][15]  (.D(values[15]), .CK(n_121_54), .Q(
      \values[65] [15]), .QN());
   DFF_X1 \values_reg[65][14]  (.D(values[14]), .CK(n_121_54), .Q(
      \values[65] [14]), .QN());
   DFF_X1 \values_reg[65][13]  (.D(values[13]), .CK(n_121_54), .Q(
      \values[65] [13]), .QN());
   DFF_X1 \values_reg[65][12]  (.D(values[12]), .CK(n_121_54), .Q(
      \values[65] [12]), .QN());
   DFF_X1 \values_reg[65][11]  (.D(values[11]), .CK(n_121_54), .Q(
      \values[65] [11]), .QN());
   DFF_X1 \values_reg[65][10]  (.D(values[10]), .CK(n_121_54), .Q(
      \values[65] [10]), .QN());
   DFF_X1 \values_reg[65][9]  (.D(values[9]), .CK(n_121_54), .Q(\values[65] [9]), 
      .QN());
   DFF_X1 \values_reg[65][8]  (.D(values[8]), .CK(n_121_54), .Q(\values[65] [8]), 
      .QN());
   DFF_X1 \values_reg[65][7]  (.D(values[7]), .CK(n_121_54), .Q(\values[65] [7]), 
      .QN());
   DFF_X1 \values_reg[65][6]  (.D(values[6]), .CK(n_121_54), .Q(\values[65] [6]), 
      .QN());
   DFF_X1 \values_reg[65][5]  (.D(values[5]), .CK(n_121_54), .Q(\values[65] [5]), 
      .QN());
   DFF_X1 \values_reg[65][4]  (.D(values[4]), .CK(n_121_54), .Q(\values[65] [4]), 
      .QN());
   DFF_X1 \values_reg[65][3]  (.D(values[3]), .CK(n_121_54), .Q(\values[65] [3]), 
      .QN());
   DFF_X1 \values_reg[65][2]  (.D(values[2]), .CK(n_121_54), .Q(\values[65] [2]), 
      .QN());
   DFF_X1 \values_reg[65][1]  (.D(values[1]), .CK(n_121_54), .Q(\values[65] [1]), 
      .QN());
   DFF_X1 \values_reg[65][0]  (.D(values[0]), .CK(n_121_54), .Q(\values[65] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[64]_reg  (.CK(clk), .E(n_64), .SE(1'b0), 
      .GCK(n_121_55));
   DFF_X1 \values_reg[64][15]  (.D(values[15]), .CK(n_121_55), .Q(
      \values[64] [15]), .QN());
   DFF_X1 \values_reg[64][14]  (.D(values[14]), .CK(n_121_55), .Q(
      \values[64] [14]), .QN());
   DFF_X1 \values_reg[64][13]  (.D(values[13]), .CK(n_121_55), .Q(
      \values[64] [13]), .QN());
   DFF_X1 \values_reg[64][12]  (.D(values[12]), .CK(n_121_55), .Q(
      \values[64] [12]), .QN());
   DFF_X1 \values_reg[64][11]  (.D(values[11]), .CK(n_121_55), .Q(
      \values[64] [11]), .QN());
   DFF_X1 \values_reg[64][10]  (.D(values[10]), .CK(n_121_55), .Q(
      \values[64] [10]), .QN());
   DFF_X1 \values_reg[64][9]  (.D(values[9]), .CK(n_121_55), .Q(\values[64] [9]), 
      .QN());
   DFF_X1 \values_reg[64][8]  (.D(values[8]), .CK(n_121_55), .Q(\values[64] [8]), 
      .QN());
   DFF_X1 \values_reg[64][7]  (.D(values[7]), .CK(n_121_55), .Q(\values[64] [7]), 
      .QN());
   DFF_X1 \values_reg[64][6]  (.D(values[6]), .CK(n_121_55), .Q(\values[64] [6]), 
      .QN());
   DFF_X1 \values_reg[64][5]  (.D(values[5]), .CK(n_121_55), .Q(\values[64] [5]), 
      .QN());
   DFF_X1 \values_reg[64][4]  (.D(values[4]), .CK(n_121_55), .Q(\values[64] [4]), 
      .QN());
   DFF_X1 \values_reg[64][3]  (.D(values[3]), .CK(n_121_55), .Q(\values[64] [3]), 
      .QN());
   DFF_X1 \values_reg[64][2]  (.D(values[2]), .CK(n_121_55), .Q(\values[64] [2]), 
      .QN());
   DFF_X1 \values_reg[64][1]  (.D(values[1]), .CK(n_121_55), .Q(\values[64] [1]), 
      .QN());
   DFF_X1 \values_reg[64][0]  (.D(values[0]), .CK(n_121_55), .Q(\values[64] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[63]_reg  (.CK(clk), .E(n_63), .SE(1'b0), 
      .GCK(n_121_56));
   DFF_X1 \values_reg[63][15]  (.D(values[15]), .CK(n_121_56), .Q(
      \values[63] [15]), .QN());
   DFF_X1 \values_reg[63][14]  (.D(values[14]), .CK(n_121_56), .Q(
      \values[63] [14]), .QN());
   DFF_X1 \values_reg[63][13]  (.D(values[13]), .CK(n_121_56), .Q(
      \values[63] [13]), .QN());
   DFF_X1 \values_reg[63][12]  (.D(values[12]), .CK(n_121_56), .Q(
      \values[63] [12]), .QN());
   DFF_X1 \values_reg[63][11]  (.D(values[11]), .CK(n_121_56), .Q(
      \values[63] [11]), .QN());
   DFF_X1 \values_reg[63][10]  (.D(values[10]), .CK(n_121_56), .Q(
      \values[63] [10]), .QN());
   DFF_X1 \values_reg[63][9]  (.D(values[9]), .CK(n_121_56), .Q(\values[63] [9]), 
      .QN());
   DFF_X1 \values_reg[63][8]  (.D(values[8]), .CK(n_121_56), .Q(\values[63] [8]), 
      .QN());
   DFF_X1 \values_reg[63][7]  (.D(values[7]), .CK(n_121_56), .Q(\values[63] [7]), 
      .QN());
   DFF_X1 \values_reg[63][6]  (.D(values[6]), .CK(n_121_56), .Q(\values[63] [6]), 
      .QN());
   DFF_X1 \values_reg[63][5]  (.D(values[5]), .CK(n_121_56), .Q(\values[63] [5]), 
      .QN());
   DFF_X1 \values_reg[63][4]  (.D(values[4]), .CK(n_121_56), .Q(\values[63] [4]), 
      .QN());
   DFF_X1 \values_reg[63][3]  (.D(values[3]), .CK(n_121_56), .Q(\values[63] [3]), 
      .QN());
   DFF_X1 \values_reg[63][2]  (.D(values[2]), .CK(n_121_56), .Q(\values[63] [2]), 
      .QN());
   DFF_X1 \values_reg[63][1]  (.D(values[1]), .CK(n_121_56), .Q(\values[63] [1]), 
      .QN());
   DFF_X1 \values_reg[63][0]  (.D(values[0]), .CK(n_121_56), .Q(\values[63] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[62]_reg  (.CK(clk), .E(n_62), .SE(1'b0), 
      .GCK(n_121_57));
   DFF_X1 \values_reg[62][15]  (.D(values[15]), .CK(n_121_57), .Q(
      \values[62] [15]), .QN());
   DFF_X1 \values_reg[62][14]  (.D(values[14]), .CK(n_121_57), .Q(
      \values[62] [14]), .QN());
   DFF_X1 \values_reg[62][13]  (.D(values[13]), .CK(n_121_57), .Q(
      \values[62] [13]), .QN());
   DFF_X1 \values_reg[62][12]  (.D(values[12]), .CK(n_121_57), .Q(
      \values[62] [12]), .QN());
   DFF_X1 \values_reg[62][11]  (.D(values[11]), .CK(n_121_57), .Q(
      \values[62] [11]), .QN());
   DFF_X1 \values_reg[62][10]  (.D(values[10]), .CK(n_121_57), .Q(
      \values[62] [10]), .QN());
   DFF_X1 \values_reg[62][9]  (.D(values[9]), .CK(n_121_57), .Q(\values[62] [9]), 
      .QN());
   DFF_X1 \values_reg[62][8]  (.D(values[8]), .CK(n_121_57), .Q(\values[62] [8]), 
      .QN());
   DFF_X1 \values_reg[62][7]  (.D(values[7]), .CK(n_121_57), .Q(\values[62] [7]), 
      .QN());
   DFF_X1 \values_reg[62][6]  (.D(values[6]), .CK(n_121_57), .Q(\values[62] [6]), 
      .QN());
   DFF_X1 \values_reg[62][5]  (.D(values[5]), .CK(n_121_57), .Q(\values[62] [5]), 
      .QN());
   DFF_X1 \values_reg[62][4]  (.D(values[4]), .CK(n_121_57), .Q(\values[62] [4]), 
      .QN());
   DFF_X1 \values_reg[62][3]  (.D(values[3]), .CK(n_121_57), .Q(\values[62] [3]), 
      .QN());
   DFF_X1 \values_reg[62][2]  (.D(values[2]), .CK(n_121_57), .Q(\values[62] [2]), 
      .QN());
   DFF_X1 \values_reg[62][1]  (.D(values[1]), .CK(n_121_57), .Q(\values[62] [1]), 
      .QN());
   DFF_X1 \values_reg[62][0]  (.D(values[0]), .CK(n_121_57), .Q(\values[62] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[61]_reg  (.CK(clk), .E(n_61), .SE(1'b0), 
      .GCK(n_121_58));
   DFF_X1 \values_reg[61][15]  (.D(values[15]), .CK(n_121_58), .Q(
      \values[61] [15]), .QN());
   DFF_X1 \values_reg[61][14]  (.D(values[14]), .CK(n_121_58), .Q(
      \values[61] [14]), .QN());
   DFF_X1 \values_reg[61][13]  (.D(values[13]), .CK(n_121_58), .Q(
      \values[61] [13]), .QN());
   DFF_X1 \values_reg[61][12]  (.D(values[12]), .CK(n_121_58), .Q(
      \values[61] [12]), .QN());
   DFF_X1 \values_reg[61][11]  (.D(values[11]), .CK(n_121_58), .Q(
      \values[61] [11]), .QN());
   DFF_X1 \values_reg[61][10]  (.D(values[10]), .CK(n_121_58), .Q(
      \values[61] [10]), .QN());
   DFF_X1 \values_reg[61][9]  (.D(values[9]), .CK(n_121_58), .Q(\values[61] [9]), 
      .QN());
   DFF_X1 \values_reg[61][8]  (.D(values[8]), .CK(n_121_58), .Q(\values[61] [8]), 
      .QN());
   DFF_X1 \values_reg[61][7]  (.D(values[7]), .CK(n_121_58), .Q(\values[61] [7]), 
      .QN());
   DFF_X1 \values_reg[61][6]  (.D(values[6]), .CK(n_121_58), .Q(\values[61] [6]), 
      .QN());
   DFF_X1 \values_reg[61][5]  (.D(values[5]), .CK(n_121_58), .Q(\values[61] [5]), 
      .QN());
   DFF_X1 \values_reg[61][4]  (.D(values[4]), .CK(n_121_58), .Q(\values[61] [4]), 
      .QN());
   DFF_X1 \values_reg[61][3]  (.D(values[3]), .CK(n_121_58), .Q(\values[61] [3]), 
      .QN());
   DFF_X1 \values_reg[61][2]  (.D(values[2]), .CK(n_121_58), .Q(\values[61] [2]), 
      .QN());
   DFF_X1 \values_reg[61][1]  (.D(values[1]), .CK(n_121_58), .Q(\values[61] [1]), 
      .QN());
   DFF_X1 \values_reg[61][0]  (.D(values[0]), .CK(n_121_58), .Q(\values[61] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[60]_reg  (.CK(clk), .E(n_60), .SE(1'b0), 
      .GCK(n_121_59));
   DFF_X1 \values_reg[60][15]  (.D(values[15]), .CK(n_121_59), .Q(
      \values[60] [15]), .QN());
   DFF_X1 \values_reg[60][14]  (.D(values[14]), .CK(n_121_59), .Q(
      \values[60] [14]), .QN());
   DFF_X1 \values_reg[60][13]  (.D(values[13]), .CK(n_121_59), .Q(
      \values[60] [13]), .QN());
   DFF_X1 \values_reg[60][12]  (.D(values[12]), .CK(n_121_59), .Q(
      \values[60] [12]), .QN());
   DFF_X1 \values_reg[60][11]  (.D(values[11]), .CK(n_121_59), .Q(
      \values[60] [11]), .QN());
   DFF_X1 \values_reg[60][10]  (.D(values[10]), .CK(n_121_59), .Q(
      \values[60] [10]), .QN());
   DFF_X1 \values_reg[60][9]  (.D(values[9]), .CK(n_121_59), .Q(\values[60] [9]), 
      .QN());
   DFF_X1 \values_reg[60][8]  (.D(values[8]), .CK(n_121_59), .Q(\values[60] [8]), 
      .QN());
   DFF_X1 \values_reg[60][7]  (.D(values[7]), .CK(n_121_59), .Q(\values[60] [7]), 
      .QN());
   DFF_X1 \values_reg[60][6]  (.D(values[6]), .CK(n_121_59), .Q(\values[60] [6]), 
      .QN());
   DFF_X1 \values_reg[60][5]  (.D(values[5]), .CK(n_121_59), .Q(\values[60] [5]), 
      .QN());
   DFF_X1 \values_reg[60][4]  (.D(values[4]), .CK(n_121_59), .Q(\values[60] [4]), 
      .QN());
   DFF_X1 \values_reg[60][3]  (.D(values[3]), .CK(n_121_59), .Q(\values[60] [3]), 
      .QN());
   DFF_X1 \values_reg[60][2]  (.D(values[2]), .CK(n_121_59), .Q(\values[60] [2]), 
      .QN());
   DFF_X1 \values_reg[60][1]  (.D(values[1]), .CK(n_121_59), .Q(\values[60] [1]), 
      .QN());
   DFF_X1 \values_reg[60][0]  (.D(values[0]), .CK(n_121_59), .Q(\values[60] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[59]_reg  (.CK(clk), .E(n_59), .SE(1'b0), 
      .GCK(n_121_60));
   DFF_X1 \values_reg[59][15]  (.D(values[15]), .CK(n_121_60), .Q(
      \values[59] [15]), .QN());
   DFF_X1 \values_reg[59][14]  (.D(values[14]), .CK(n_121_60), .Q(
      \values[59] [14]), .QN());
   DFF_X1 \values_reg[59][13]  (.D(values[13]), .CK(n_121_60), .Q(
      \values[59] [13]), .QN());
   DFF_X1 \values_reg[59][12]  (.D(values[12]), .CK(n_121_60), .Q(
      \values[59] [12]), .QN());
   DFF_X1 \values_reg[59][11]  (.D(values[11]), .CK(n_121_60), .Q(
      \values[59] [11]), .QN());
   DFF_X1 \values_reg[59][10]  (.D(values[10]), .CK(n_121_60), .Q(
      \values[59] [10]), .QN());
   DFF_X1 \values_reg[59][9]  (.D(values[9]), .CK(n_121_60), .Q(\values[59] [9]), 
      .QN());
   DFF_X1 \values_reg[59][8]  (.D(values[8]), .CK(n_121_60), .Q(\values[59] [8]), 
      .QN());
   DFF_X1 \values_reg[59][7]  (.D(values[7]), .CK(n_121_60), .Q(\values[59] [7]), 
      .QN());
   DFF_X1 \values_reg[59][6]  (.D(values[6]), .CK(n_121_60), .Q(\values[59] [6]), 
      .QN());
   DFF_X1 \values_reg[59][5]  (.D(values[5]), .CK(n_121_60), .Q(\values[59] [5]), 
      .QN());
   DFF_X1 \values_reg[59][4]  (.D(values[4]), .CK(n_121_60), .Q(\values[59] [4]), 
      .QN());
   DFF_X1 \values_reg[59][3]  (.D(values[3]), .CK(n_121_60), .Q(\values[59] [3]), 
      .QN());
   DFF_X1 \values_reg[59][2]  (.D(values[2]), .CK(n_121_60), .Q(\values[59] [2]), 
      .QN());
   DFF_X1 \values_reg[59][1]  (.D(values[1]), .CK(n_121_60), .Q(\values[59] [1]), 
      .QN());
   DFF_X1 \values_reg[59][0]  (.D(values[0]), .CK(n_121_60), .Q(\values[59] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[58]_reg  (.CK(clk), .E(n_58), .SE(1'b0), 
      .GCK(n_121_61));
   DFF_X1 \values_reg[58][15]  (.D(values[15]), .CK(n_121_61), .Q(
      \values[58] [15]), .QN());
   DFF_X1 \values_reg[58][14]  (.D(values[14]), .CK(n_121_61), .Q(
      \values[58] [14]), .QN());
   DFF_X1 \values_reg[58][13]  (.D(values[13]), .CK(n_121_61), .Q(
      \values[58] [13]), .QN());
   DFF_X1 \values_reg[58][12]  (.D(values[12]), .CK(n_121_61), .Q(
      \values[58] [12]), .QN());
   DFF_X1 \values_reg[58][11]  (.D(values[11]), .CK(n_121_61), .Q(
      \values[58] [11]), .QN());
   DFF_X1 \values_reg[58][10]  (.D(values[10]), .CK(n_121_61), .Q(
      \values[58] [10]), .QN());
   DFF_X1 \values_reg[58][9]  (.D(values[9]), .CK(n_121_61), .Q(\values[58] [9]), 
      .QN());
   DFF_X1 \values_reg[58][8]  (.D(values[8]), .CK(n_121_61), .Q(\values[58] [8]), 
      .QN());
   DFF_X1 \values_reg[58][7]  (.D(values[7]), .CK(n_121_61), .Q(\values[58] [7]), 
      .QN());
   DFF_X1 \values_reg[58][6]  (.D(values[6]), .CK(n_121_61), .Q(\values[58] [6]), 
      .QN());
   DFF_X1 \values_reg[58][5]  (.D(values[5]), .CK(n_121_61), .Q(\values[58] [5]), 
      .QN());
   DFF_X1 \values_reg[58][4]  (.D(values[4]), .CK(n_121_61), .Q(\values[58] [4]), 
      .QN());
   DFF_X1 \values_reg[58][3]  (.D(values[3]), .CK(n_121_61), .Q(\values[58] [3]), 
      .QN());
   DFF_X1 \values_reg[58][2]  (.D(values[2]), .CK(n_121_61), .Q(\values[58] [2]), 
      .QN());
   DFF_X1 \values_reg[58][1]  (.D(values[1]), .CK(n_121_61), .Q(\values[58] [1]), 
      .QN());
   DFF_X1 \values_reg[58][0]  (.D(values[0]), .CK(n_121_61), .Q(\values[58] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[57]_reg  (.CK(clk), .E(n_57), .SE(1'b0), 
      .GCK(n_121_62));
   DFF_X1 \values_reg[57][15]  (.D(values[15]), .CK(n_121_62), .Q(
      \values[57] [15]), .QN());
   DFF_X1 \values_reg[57][14]  (.D(values[14]), .CK(n_121_62), .Q(
      \values[57] [14]), .QN());
   DFF_X1 \values_reg[57][13]  (.D(values[13]), .CK(n_121_62), .Q(
      \values[57] [13]), .QN());
   DFF_X1 \values_reg[57][12]  (.D(values[12]), .CK(n_121_62), .Q(
      \values[57] [12]), .QN());
   DFF_X1 \values_reg[57][11]  (.D(values[11]), .CK(n_121_62), .Q(
      \values[57] [11]), .QN());
   DFF_X1 \values_reg[57][10]  (.D(values[10]), .CK(n_121_62), .Q(
      \values[57] [10]), .QN());
   DFF_X1 \values_reg[57][9]  (.D(values[9]), .CK(n_121_62), .Q(\values[57] [9]), 
      .QN());
   DFF_X1 \values_reg[57][8]  (.D(values[8]), .CK(n_121_62), .Q(\values[57] [8]), 
      .QN());
   DFF_X1 \values_reg[57][7]  (.D(values[7]), .CK(n_121_62), .Q(\values[57] [7]), 
      .QN());
   DFF_X1 \values_reg[57][6]  (.D(values[6]), .CK(n_121_62), .Q(\values[57] [6]), 
      .QN());
   DFF_X1 \values_reg[57][5]  (.D(values[5]), .CK(n_121_62), .Q(\values[57] [5]), 
      .QN());
   DFF_X1 \values_reg[57][4]  (.D(values[4]), .CK(n_121_62), .Q(\values[57] [4]), 
      .QN());
   DFF_X1 \values_reg[57][3]  (.D(values[3]), .CK(n_121_62), .Q(\values[57] [3]), 
      .QN());
   DFF_X1 \values_reg[57][2]  (.D(values[2]), .CK(n_121_62), .Q(\values[57] [2]), 
      .QN());
   DFF_X1 \values_reg[57][1]  (.D(values[1]), .CK(n_121_62), .Q(\values[57] [1]), 
      .QN());
   DFF_X1 \values_reg[57][0]  (.D(values[0]), .CK(n_121_62), .Q(\values[57] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[56]_reg  (.CK(clk), .E(n_56), .SE(1'b0), 
      .GCK(n_121_63));
   DFF_X1 \values_reg[56][15]  (.D(values[15]), .CK(n_121_63), .Q(
      \values[56] [15]), .QN());
   DFF_X1 \values_reg[56][14]  (.D(values[14]), .CK(n_121_63), .Q(
      \values[56] [14]), .QN());
   DFF_X1 \values_reg[56][13]  (.D(values[13]), .CK(n_121_63), .Q(
      \values[56] [13]), .QN());
   DFF_X1 \values_reg[56][12]  (.D(values[12]), .CK(n_121_63), .Q(
      \values[56] [12]), .QN());
   DFF_X1 \values_reg[56][11]  (.D(values[11]), .CK(n_121_63), .Q(
      \values[56] [11]), .QN());
   DFF_X1 \values_reg[56][10]  (.D(values[10]), .CK(n_121_63), .Q(
      \values[56] [10]), .QN());
   DFF_X1 \values_reg[56][9]  (.D(values[9]), .CK(n_121_63), .Q(\values[56] [9]), 
      .QN());
   DFF_X1 \values_reg[56][8]  (.D(values[8]), .CK(n_121_63), .Q(\values[56] [8]), 
      .QN());
   DFF_X1 \values_reg[56][7]  (.D(values[7]), .CK(n_121_63), .Q(\values[56] [7]), 
      .QN());
   DFF_X1 \values_reg[56][6]  (.D(values[6]), .CK(n_121_63), .Q(\values[56] [6]), 
      .QN());
   DFF_X1 \values_reg[56][5]  (.D(values[5]), .CK(n_121_63), .Q(\values[56] [5]), 
      .QN());
   DFF_X1 \values_reg[56][4]  (.D(values[4]), .CK(n_121_63), .Q(\values[56] [4]), 
      .QN());
   DFF_X1 \values_reg[56][3]  (.D(values[3]), .CK(n_121_63), .Q(\values[56] [3]), 
      .QN());
   DFF_X1 \values_reg[56][2]  (.D(values[2]), .CK(n_121_63), .Q(\values[56] [2]), 
      .QN());
   DFF_X1 \values_reg[56][1]  (.D(values[1]), .CK(n_121_63), .Q(\values[56] [1]), 
      .QN());
   DFF_X1 \values_reg[56][0]  (.D(values[0]), .CK(n_121_63), .Q(\values[56] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[55]_reg  (.CK(clk), .E(n_55), .SE(1'b0), 
      .GCK(n_121_64));
   DFF_X1 \values_reg[55][15]  (.D(values[15]), .CK(n_121_64), .Q(
      \values[55] [15]), .QN());
   DFF_X1 \values_reg[55][14]  (.D(values[14]), .CK(n_121_64), .Q(
      \values[55] [14]), .QN());
   DFF_X1 \values_reg[55][13]  (.D(values[13]), .CK(n_121_64), .Q(
      \values[55] [13]), .QN());
   DFF_X1 \values_reg[55][12]  (.D(values[12]), .CK(n_121_64), .Q(
      \values[55] [12]), .QN());
   DFF_X1 \values_reg[55][11]  (.D(values[11]), .CK(n_121_64), .Q(
      \values[55] [11]), .QN());
   DFF_X1 \values_reg[55][10]  (.D(values[10]), .CK(n_121_64), .Q(
      \values[55] [10]), .QN());
   DFF_X1 \values_reg[55][9]  (.D(values[9]), .CK(n_121_64), .Q(\values[55] [9]), 
      .QN());
   DFF_X1 \values_reg[55][8]  (.D(values[8]), .CK(n_121_64), .Q(\values[55] [8]), 
      .QN());
   DFF_X1 \values_reg[55][7]  (.D(values[7]), .CK(n_121_64), .Q(\values[55] [7]), 
      .QN());
   DFF_X1 \values_reg[55][6]  (.D(values[6]), .CK(n_121_64), .Q(\values[55] [6]), 
      .QN());
   DFF_X1 \values_reg[55][5]  (.D(values[5]), .CK(n_121_64), .Q(\values[55] [5]), 
      .QN());
   DFF_X1 \values_reg[55][4]  (.D(values[4]), .CK(n_121_64), .Q(\values[55] [4]), 
      .QN());
   DFF_X1 \values_reg[55][3]  (.D(values[3]), .CK(n_121_64), .Q(\values[55] [3]), 
      .QN());
   DFF_X1 \values_reg[55][2]  (.D(values[2]), .CK(n_121_64), .Q(\values[55] [2]), 
      .QN());
   DFF_X1 \values_reg[55][1]  (.D(values[1]), .CK(n_121_64), .Q(\values[55] [1]), 
      .QN());
   DFF_X1 \values_reg[55][0]  (.D(values[0]), .CK(n_121_64), .Q(\values[55] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[54]_reg  (.CK(clk), .E(n_54), .SE(1'b0), 
      .GCK(n_121_65));
   DFF_X1 \values_reg[54][15]  (.D(values[15]), .CK(n_121_65), .Q(
      \values[54] [15]), .QN());
   DFF_X1 \values_reg[54][14]  (.D(values[14]), .CK(n_121_65), .Q(
      \values[54] [14]), .QN());
   DFF_X1 \values_reg[54][13]  (.D(values[13]), .CK(n_121_65), .Q(
      \values[54] [13]), .QN());
   DFF_X1 \values_reg[54][12]  (.D(values[12]), .CK(n_121_65), .Q(
      \values[54] [12]), .QN());
   DFF_X1 \values_reg[54][11]  (.D(values[11]), .CK(n_121_65), .Q(
      \values[54] [11]), .QN());
   DFF_X1 \values_reg[54][10]  (.D(values[10]), .CK(n_121_65), .Q(
      \values[54] [10]), .QN());
   DFF_X1 \values_reg[54][9]  (.D(values[9]), .CK(n_121_65), .Q(\values[54] [9]), 
      .QN());
   DFF_X1 \values_reg[54][8]  (.D(values[8]), .CK(n_121_65), .Q(\values[54] [8]), 
      .QN());
   DFF_X1 \values_reg[54][7]  (.D(values[7]), .CK(n_121_65), .Q(\values[54] [7]), 
      .QN());
   DFF_X1 \values_reg[54][6]  (.D(values[6]), .CK(n_121_65), .Q(\values[54] [6]), 
      .QN());
   DFF_X1 \values_reg[54][5]  (.D(values[5]), .CK(n_121_65), .Q(\values[54] [5]), 
      .QN());
   DFF_X1 \values_reg[54][4]  (.D(values[4]), .CK(n_121_65), .Q(\values[54] [4]), 
      .QN());
   DFF_X1 \values_reg[54][3]  (.D(values[3]), .CK(n_121_65), .Q(\values[54] [3]), 
      .QN());
   DFF_X1 \values_reg[54][2]  (.D(values[2]), .CK(n_121_65), .Q(\values[54] [2]), 
      .QN());
   DFF_X1 \values_reg[54][1]  (.D(values[1]), .CK(n_121_65), .Q(\values[54] [1]), 
      .QN());
   DFF_X1 \values_reg[54][0]  (.D(values[0]), .CK(n_121_65), .Q(\values[54] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[53]_reg  (.CK(clk), .E(n_53), .SE(1'b0), 
      .GCK(n_121_66));
   DFF_X1 \values_reg[53][15]  (.D(values[15]), .CK(n_121_66), .Q(
      \values[53] [15]), .QN());
   DFF_X1 \values_reg[53][14]  (.D(values[14]), .CK(n_121_66), .Q(
      \values[53] [14]), .QN());
   DFF_X1 \values_reg[53][13]  (.D(values[13]), .CK(n_121_66), .Q(
      \values[53] [13]), .QN());
   DFF_X1 \values_reg[53][12]  (.D(values[12]), .CK(n_121_66), .Q(
      \values[53] [12]), .QN());
   DFF_X1 \values_reg[53][11]  (.D(values[11]), .CK(n_121_66), .Q(
      \values[53] [11]), .QN());
   DFF_X1 \values_reg[53][10]  (.D(values[10]), .CK(n_121_66), .Q(
      \values[53] [10]), .QN());
   DFF_X1 \values_reg[53][9]  (.D(values[9]), .CK(n_121_66), .Q(\values[53] [9]), 
      .QN());
   DFF_X1 \values_reg[53][8]  (.D(values[8]), .CK(n_121_66), .Q(\values[53] [8]), 
      .QN());
   DFF_X1 \values_reg[53][7]  (.D(values[7]), .CK(n_121_66), .Q(\values[53] [7]), 
      .QN());
   DFF_X1 \values_reg[53][6]  (.D(values[6]), .CK(n_121_66), .Q(\values[53] [6]), 
      .QN());
   DFF_X1 \values_reg[53][5]  (.D(values[5]), .CK(n_121_66), .Q(\values[53] [5]), 
      .QN());
   DFF_X1 \values_reg[53][4]  (.D(values[4]), .CK(n_121_66), .Q(\values[53] [4]), 
      .QN());
   DFF_X1 \values_reg[53][3]  (.D(values[3]), .CK(n_121_66), .Q(\values[53] [3]), 
      .QN());
   DFF_X1 \values_reg[53][2]  (.D(values[2]), .CK(n_121_66), .Q(\values[53] [2]), 
      .QN());
   DFF_X1 \values_reg[53][1]  (.D(values[1]), .CK(n_121_66), .Q(\values[53] [1]), 
      .QN());
   DFF_X1 \values_reg[53][0]  (.D(values[0]), .CK(n_121_66), .Q(\values[53] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[52]_reg  (.CK(clk), .E(n_52), .SE(1'b0), 
      .GCK(n_121_67));
   DFF_X1 \values_reg[52][15]  (.D(values[15]), .CK(n_121_67), .Q(
      \values[52] [15]), .QN());
   DFF_X1 \values_reg[52][14]  (.D(values[14]), .CK(n_121_67), .Q(
      \values[52] [14]), .QN());
   DFF_X1 \values_reg[52][13]  (.D(values[13]), .CK(n_121_67), .Q(
      \values[52] [13]), .QN());
   DFF_X1 \values_reg[52][12]  (.D(values[12]), .CK(n_121_67), .Q(
      \values[52] [12]), .QN());
   DFF_X1 \values_reg[52][11]  (.D(values[11]), .CK(n_121_67), .Q(
      \values[52] [11]), .QN());
   DFF_X1 \values_reg[52][10]  (.D(values[10]), .CK(n_121_67), .Q(
      \values[52] [10]), .QN());
   DFF_X1 \values_reg[52][9]  (.D(values[9]), .CK(n_121_67), .Q(\values[52] [9]), 
      .QN());
   DFF_X1 \values_reg[52][8]  (.D(values[8]), .CK(n_121_67), .Q(\values[52] [8]), 
      .QN());
   DFF_X1 \values_reg[52][7]  (.D(values[7]), .CK(n_121_67), .Q(\values[52] [7]), 
      .QN());
   DFF_X1 \values_reg[52][6]  (.D(values[6]), .CK(n_121_67), .Q(\values[52] [6]), 
      .QN());
   DFF_X1 \values_reg[52][5]  (.D(values[5]), .CK(n_121_67), .Q(\values[52] [5]), 
      .QN());
   DFF_X1 \values_reg[52][4]  (.D(values[4]), .CK(n_121_67), .Q(\values[52] [4]), 
      .QN());
   DFF_X1 \values_reg[52][3]  (.D(values[3]), .CK(n_121_67), .Q(\values[52] [3]), 
      .QN());
   DFF_X1 \values_reg[52][2]  (.D(values[2]), .CK(n_121_67), .Q(\values[52] [2]), 
      .QN());
   DFF_X1 \values_reg[52][1]  (.D(values[1]), .CK(n_121_67), .Q(\values[52] [1]), 
      .QN());
   DFF_X1 \values_reg[52][0]  (.D(values[0]), .CK(n_121_67), .Q(\values[52] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[51]_reg  (.CK(clk), .E(n_51), .SE(1'b0), 
      .GCK(n_121_68));
   DFF_X1 \values_reg[51][15]  (.D(values[15]), .CK(n_121_68), .Q(
      \values[51] [15]), .QN());
   DFF_X1 \values_reg[51][14]  (.D(values[14]), .CK(n_121_68), .Q(
      \values[51] [14]), .QN());
   DFF_X1 \values_reg[51][13]  (.D(values[13]), .CK(n_121_68), .Q(
      \values[51] [13]), .QN());
   DFF_X1 \values_reg[51][12]  (.D(values[12]), .CK(n_121_68), .Q(
      \values[51] [12]), .QN());
   DFF_X1 \values_reg[51][11]  (.D(values[11]), .CK(n_121_68), .Q(
      \values[51] [11]), .QN());
   DFF_X1 \values_reg[51][10]  (.D(values[10]), .CK(n_121_68), .Q(
      \values[51] [10]), .QN());
   DFF_X1 \values_reg[51][9]  (.D(values[9]), .CK(n_121_68), .Q(\values[51] [9]), 
      .QN());
   DFF_X1 \values_reg[51][8]  (.D(values[8]), .CK(n_121_68), .Q(\values[51] [8]), 
      .QN());
   DFF_X1 \values_reg[51][7]  (.D(values[7]), .CK(n_121_68), .Q(\values[51] [7]), 
      .QN());
   DFF_X1 \values_reg[51][6]  (.D(values[6]), .CK(n_121_68), .Q(\values[51] [6]), 
      .QN());
   DFF_X1 \values_reg[51][5]  (.D(values[5]), .CK(n_121_68), .Q(\values[51] [5]), 
      .QN());
   DFF_X1 \values_reg[51][4]  (.D(values[4]), .CK(n_121_68), .Q(\values[51] [4]), 
      .QN());
   DFF_X1 \values_reg[51][3]  (.D(values[3]), .CK(n_121_68), .Q(\values[51] [3]), 
      .QN());
   DFF_X1 \values_reg[51][2]  (.D(values[2]), .CK(n_121_68), .Q(\values[51] [2]), 
      .QN());
   DFF_X1 \values_reg[51][1]  (.D(values[1]), .CK(n_121_68), .Q(\values[51] [1]), 
      .QN());
   DFF_X1 \values_reg[51][0]  (.D(values[0]), .CK(n_121_68), .Q(\values[51] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[50]_reg  (.CK(clk), .E(n_50), .SE(1'b0), 
      .GCK(n_121_69));
   DFF_X1 \values_reg[50][15]  (.D(values[15]), .CK(n_121_69), .Q(
      \values[50] [15]), .QN());
   DFF_X1 \values_reg[50][14]  (.D(values[14]), .CK(n_121_69), .Q(
      \values[50] [14]), .QN());
   DFF_X1 \values_reg[50][13]  (.D(values[13]), .CK(n_121_69), .Q(
      \values[50] [13]), .QN());
   DFF_X1 \values_reg[50][12]  (.D(values[12]), .CK(n_121_69), .Q(
      \values[50] [12]), .QN());
   DFF_X1 \values_reg[50][11]  (.D(values[11]), .CK(n_121_69), .Q(
      \values[50] [11]), .QN());
   DFF_X1 \values_reg[50][10]  (.D(values[10]), .CK(n_121_69), .Q(
      \values[50] [10]), .QN());
   DFF_X1 \values_reg[50][9]  (.D(values[9]), .CK(n_121_69), .Q(\values[50] [9]), 
      .QN());
   DFF_X1 \values_reg[50][8]  (.D(values[8]), .CK(n_121_69), .Q(\values[50] [8]), 
      .QN());
   DFF_X1 \values_reg[50][7]  (.D(values[7]), .CK(n_121_69), .Q(\values[50] [7]), 
      .QN());
   DFF_X1 \values_reg[50][6]  (.D(values[6]), .CK(n_121_69), .Q(\values[50] [6]), 
      .QN());
   DFF_X1 \values_reg[50][5]  (.D(values[5]), .CK(n_121_69), .Q(\values[50] [5]), 
      .QN());
   DFF_X1 \values_reg[50][4]  (.D(values[4]), .CK(n_121_69), .Q(\values[50] [4]), 
      .QN());
   DFF_X1 \values_reg[50][3]  (.D(values[3]), .CK(n_121_69), .Q(\values[50] [3]), 
      .QN());
   DFF_X1 \values_reg[50][2]  (.D(values[2]), .CK(n_121_69), .Q(\values[50] [2]), 
      .QN());
   DFF_X1 \values_reg[50][1]  (.D(values[1]), .CK(n_121_69), .Q(\values[50] [1]), 
      .QN());
   DFF_X1 \values_reg[50][0]  (.D(values[0]), .CK(n_121_69), .Q(\values[50] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[49]_reg  (.CK(clk), .E(n_49), .SE(1'b0), 
      .GCK(n_121_70));
   DFF_X1 \values_reg[49][15]  (.D(values[15]), .CK(n_121_70), .Q(
      \values[49] [15]), .QN());
   DFF_X1 \values_reg[49][14]  (.D(values[14]), .CK(n_121_70), .Q(
      \values[49] [14]), .QN());
   DFF_X1 \values_reg[49][13]  (.D(values[13]), .CK(n_121_70), .Q(
      \values[49] [13]), .QN());
   DFF_X1 \values_reg[49][12]  (.D(values[12]), .CK(n_121_70), .Q(
      \values[49] [12]), .QN());
   DFF_X1 \values_reg[49][11]  (.D(values[11]), .CK(n_121_70), .Q(
      \values[49] [11]), .QN());
   DFF_X1 \values_reg[49][10]  (.D(values[10]), .CK(n_121_70), .Q(
      \values[49] [10]), .QN());
   DFF_X1 \values_reg[49][9]  (.D(values[9]), .CK(n_121_70), .Q(\values[49] [9]), 
      .QN());
   DFF_X1 \values_reg[49][8]  (.D(values[8]), .CK(n_121_70), .Q(\values[49] [8]), 
      .QN());
   DFF_X1 \values_reg[49][7]  (.D(values[7]), .CK(n_121_70), .Q(\values[49] [7]), 
      .QN());
   DFF_X1 \values_reg[49][6]  (.D(values[6]), .CK(n_121_70), .Q(\values[49] [6]), 
      .QN());
   DFF_X1 \values_reg[49][5]  (.D(values[5]), .CK(n_121_70), .Q(\values[49] [5]), 
      .QN());
   DFF_X1 \values_reg[49][4]  (.D(values[4]), .CK(n_121_70), .Q(\values[49] [4]), 
      .QN());
   DFF_X1 \values_reg[49][3]  (.D(values[3]), .CK(n_121_70), .Q(\values[49] [3]), 
      .QN());
   DFF_X1 \values_reg[49][2]  (.D(values[2]), .CK(n_121_70), .Q(\values[49] [2]), 
      .QN());
   DFF_X1 \values_reg[49][1]  (.D(values[1]), .CK(n_121_70), .Q(\values[49] [1]), 
      .QN());
   DFF_X1 \values_reg[49][0]  (.D(values[0]), .CK(n_121_70), .Q(\values[49] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[48]_reg  (.CK(clk), .E(n_48), .SE(1'b0), 
      .GCK(n_121_71));
   DFF_X1 \values_reg[48][15]  (.D(values[15]), .CK(n_121_71), .Q(
      \values[48] [15]), .QN());
   DFF_X1 \values_reg[48][14]  (.D(values[14]), .CK(n_121_71), .Q(
      \values[48] [14]), .QN());
   DFF_X1 \values_reg[48][13]  (.D(values[13]), .CK(n_121_71), .Q(
      \values[48] [13]), .QN());
   DFF_X1 \values_reg[48][12]  (.D(values[12]), .CK(n_121_71), .Q(
      \values[48] [12]), .QN());
   DFF_X1 \values_reg[48][11]  (.D(values[11]), .CK(n_121_71), .Q(
      \values[48] [11]), .QN());
   DFF_X1 \values_reg[48][10]  (.D(values[10]), .CK(n_121_71), .Q(
      \values[48] [10]), .QN());
   DFF_X1 \values_reg[48][9]  (.D(values[9]), .CK(n_121_71), .Q(\values[48] [9]), 
      .QN());
   DFF_X1 \values_reg[48][8]  (.D(values[8]), .CK(n_121_71), .Q(\values[48] [8]), 
      .QN());
   DFF_X1 \values_reg[48][7]  (.D(values[7]), .CK(n_121_71), .Q(\values[48] [7]), 
      .QN());
   DFF_X1 \values_reg[48][6]  (.D(values[6]), .CK(n_121_71), .Q(\values[48] [6]), 
      .QN());
   DFF_X1 \values_reg[48][5]  (.D(values[5]), .CK(n_121_71), .Q(\values[48] [5]), 
      .QN());
   DFF_X1 \values_reg[48][4]  (.D(values[4]), .CK(n_121_71), .Q(\values[48] [4]), 
      .QN());
   DFF_X1 \values_reg[48][3]  (.D(values[3]), .CK(n_121_71), .Q(\values[48] [3]), 
      .QN());
   DFF_X1 \values_reg[48][2]  (.D(values[2]), .CK(n_121_71), .Q(\values[48] [2]), 
      .QN());
   DFF_X1 \values_reg[48][1]  (.D(values[1]), .CK(n_121_71), .Q(\values[48] [1]), 
      .QN());
   DFF_X1 \values_reg[48][0]  (.D(values[0]), .CK(n_121_71), .Q(\values[48] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[47]_reg  (.CK(clk), .E(n_47), .SE(1'b0), 
      .GCK(n_121_72));
   DFF_X1 \values_reg[47][15]  (.D(values[15]), .CK(n_121_72), .Q(
      \values[47] [15]), .QN());
   DFF_X1 \values_reg[47][14]  (.D(values[14]), .CK(n_121_72), .Q(
      \values[47] [14]), .QN());
   DFF_X1 \values_reg[47][13]  (.D(values[13]), .CK(n_121_72), .Q(
      \values[47] [13]), .QN());
   DFF_X1 \values_reg[47][12]  (.D(values[12]), .CK(n_121_72), .Q(
      \values[47] [12]), .QN());
   DFF_X1 \values_reg[47][11]  (.D(values[11]), .CK(n_121_72), .Q(
      \values[47] [11]), .QN());
   DFF_X1 \values_reg[47][10]  (.D(values[10]), .CK(n_121_72), .Q(
      \values[47] [10]), .QN());
   DFF_X1 \values_reg[47][9]  (.D(values[9]), .CK(n_121_72), .Q(\values[47] [9]), 
      .QN());
   DFF_X1 \values_reg[47][8]  (.D(values[8]), .CK(n_121_72), .Q(\values[47] [8]), 
      .QN());
   DFF_X1 \values_reg[47][7]  (.D(values[7]), .CK(n_121_72), .Q(\values[47] [7]), 
      .QN());
   DFF_X1 \values_reg[47][6]  (.D(values[6]), .CK(n_121_72), .Q(\values[47] [6]), 
      .QN());
   DFF_X1 \values_reg[47][5]  (.D(values[5]), .CK(n_121_72), .Q(\values[47] [5]), 
      .QN());
   DFF_X1 \values_reg[47][4]  (.D(values[4]), .CK(n_121_72), .Q(\values[47] [4]), 
      .QN());
   DFF_X1 \values_reg[47][3]  (.D(values[3]), .CK(n_121_72), .Q(\values[47] [3]), 
      .QN());
   DFF_X1 \values_reg[47][2]  (.D(values[2]), .CK(n_121_72), .Q(\values[47] [2]), 
      .QN());
   DFF_X1 \values_reg[47][1]  (.D(values[1]), .CK(n_121_72), .Q(\values[47] [1]), 
      .QN());
   DFF_X1 \values_reg[47][0]  (.D(values[0]), .CK(n_121_72), .Q(\values[47] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[46]_reg  (.CK(clk), .E(n_46), .SE(1'b0), 
      .GCK(n_121_73));
   DFF_X1 \values_reg[46][15]  (.D(values[15]), .CK(n_121_73), .Q(
      \values[46] [15]), .QN());
   DFF_X1 \values_reg[46][14]  (.D(values[14]), .CK(n_121_73), .Q(
      \values[46] [14]), .QN());
   DFF_X1 \values_reg[46][13]  (.D(values[13]), .CK(n_121_73), .Q(
      \values[46] [13]), .QN());
   DFF_X1 \values_reg[46][12]  (.D(values[12]), .CK(n_121_73), .Q(
      \values[46] [12]), .QN());
   DFF_X1 \values_reg[46][11]  (.D(values[11]), .CK(n_121_73), .Q(
      \values[46] [11]), .QN());
   DFF_X1 \values_reg[46][10]  (.D(values[10]), .CK(n_121_73), .Q(
      \values[46] [10]), .QN());
   DFF_X1 \values_reg[46][9]  (.D(values[9]), .CK(n_121_73), .Q(\values[46] [9]), 
      .QN());
   DFF_X1 \values_reg[46][8]  (.D(values[8]), .CK(n_121_73), .Q(\values[46] [8]), 
      .QN());
   DFF_X1 \values_reg[46][7]  (.D(values[7]), .CK(n_121_73), .Q(\values[46] [7]), 
      .QN());
   DFF_X1 \values_reg[46][6]  (.D(values[6]), .CK(n_121_73), .Q(\values[46] [6]), 
      .QN());
   DFF_X1 \values_reg[46][5]  (.D(values[5]), .CK(n_121_73), .Q(\values[46] [5]), 
      .QN());
   DFF_X1 \values_reg[46][4]  (.D(values[4]), .CK(n_121_73), .Q(\values[46] [4]), 
      .QN());
   DFF_X1 \values_reg[46][3]  (.D(values[3]), .CK(n_121_73), .Q(\values[46] [3]), 
      .QN());
   DFF_X1 \values_reg[46][2]  (.D(values[2]), .CK(n_121_73), .Q(\values[46] [2]), 
      .QN());
   DFF_X1 \values_reg[46][1]  (.D(values[1]), .CK(n_121_73), .Q(\values[46] [1]), 
      .QN());
   DFF_X1 \values_reg[46][0]  (.D(values[0]), .CK(n_121_73), .Q(\values[46] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[45]_reg  (.CK(clk), .E(n_45), .SE(1'b0), 
      .GCK(n_121_74));
   DFF_X1 \values_reg[45][15]  (.D(values[15]), .CK(n_121_74), .Q(
      \values[45] [15]), .QN());
   DFF_X1 \values_reg[45][14]  (.D(values[14]), .CK(n_121_74), .Q(
      \values[45] [14]), .QN());
   DFF_X1 \values_reg[45][13]  (.D(values[13]), .CK(n_121_74), .Q(
      \values[45] [13]), .QN());
   DFF_X1 \values_reg[45][12]  (.D(values[12]), .CK(n_121_74), .Q(
      \values[45] [12]), .QN());
   DFF_X1 \values_reg[45][11]  (.D(values[11]), .CK(n_121_74), .Q(
      \values[45] [11]), .QN());
   DFF_X1 \values_reg[45][10]  (.D(values[10]), .CK(n_121_74), .Q(
      \values[45] [10]), .QN());
   DFF_X1 \values_reg[45][9]  (.D(values[9]), .CK(n_121_74), .Q(\values[45] [9]), 
      .QN());
   DFF_X1 \values_reg[45][8]  (.D(values[8]), .CK(n_121_74), .Q(\values[45] [8]), 
      .QN());
   DFF_X1 \values_reg[45][7]  (.D(values[7]), .CK(n_121_74), .Q(\values[45] [7]), 
      .QN());
   DFF_X1 \values_reg[45][6]  (.D(values[6]), .CK(n_121_74), .Q(\values[45] [6]), 
      .QN());
   DFF_X1 \values_reg[45][5]  (.D(values[5]), .CK(n_121_74), .Q(\values[45] [5]), 
      .QN());
   DFF_X1 \values_reg[45][4]  (.D(values[4]), .CK(n_121_74), .Q(\values[45] [4]), 
      .QN());
   DFF_X1 \values_reg[45][3]  (.D(values[3]), .CK(n_121_74), .Q(\values[45] [3]), 
      .QN());
   DFF_X1 \values_reg[45][2]  (.D(values[2]), .CK(n_121_74), .Q(\values[45] [2]), 
      .QN());
   DFF_X1 \values_reg[45][1]  (.D(values[1]), .CK(n_121_74), .Q(\values[45] [1]), 
      .QN());
   DFF_X1 \values_reg[45][0]  (.D(values[0]), .CK(n_121_74), .Q(\values[45] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[44]_reg  (.CK(clk), .E(n_44), .SE(1'b0), 
      .GCK(n_121_75));
   DFF_X1 \values_reg[44][15]  (.D(values[15]), .CK(n_121_75), .Q(
      \values[44] [15]), .QN());
   DFF_X1 \values_reg[44][14]  (.D(values[14]), .CK(n_121_75), .Q(
      \values[44] [14]), .QN());
   DFF_X1 \values_reg[44][13]  (.D(values[13]), .CK(n_121_75), .Q(
      \values[44] [13]), .QN());
   DFF_X1 \values_reg[44][12]  (.D(values[12]), .CK(n_121_75), .Q(
      \values[44] [12]), .QN());
   DFF_X1 \values_reg[44][11]  (.D(values[11]), .CK(n_121_75), .Q(
      \values[44] [11]), .QN());
   DFF_X1 \values_reg[44][10]  (.D(values[10]), .CK(n_121_75), .Q(
      \values[44] [10]), .QN());
   DFF_X1 \values_reg[44][9]  (.D(values[9]), .CK(n_121_75), .Q(\values[44] [9]), 
      .QN());
   DFF_X1 \values_reg[44][8]  (.D(values[8]), .CK(n_121_75), .Q(\values[44] [8]), 
      .QN());
   DFF_X1 \values_reg[44][7]  (.D(values[7]), .CK(n_121_75), .Q(\values[44] [7]), 
      .QN());
   DFF_X1 \values_reg[44][6]  (.D(values[6]), .CK(n_121_75), .Q(\values[44] [6]), 
      .QN());
   DFF_X1 \values_reg[44][5]  (.D(values[5]), .CK(n_121_75), .Q(\values[44] [5]), 
      .QN());
   DFF_X1 \values_reg[44][4]  (.D(values[4]), .CK(n_121_75), .Q(\values[44] [4]), 
      .QN());
   DFF_X1 \values_reg[44][3]  (.D(values[3]), .CK(n_121_75), .Q(\values[44] [3]), 
      .QN());
   DFF_X1 \values_reg[44][2]  (.D(values[2]), .CK(n_121_75), .Q(\values[44] [2]), 
      .QN());
   DFF_X1 \values_reg[44][1]  (.D(values[1]), .CK(n_121_75), .Q(\values[44] [1]), 
      .QN());
   DFF_X1 \values_reg[44][0]  (.D(values[0]), .CK(n_121_75), .Q(\values[44] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[43]_reg  (.CK(clk), .E(n_43), .SE(1'b0), 
      .GCK(n_121_76));
   DFF_X1 \values_reg[43][15]  (.D(values[15]), .CK(n_121_76), .Q(
      \values[43] [15]), .QN());
   DFF_X1 \values_reg[43][14]  (.D(values[14]), .CK(n_121_76), .Q(
      \values[43] [14]), .QN());
   DFF_X1 \values_reg[43][13]  (.D(values[13]), .CK(n_121_76), .Q(
      \values[43] [13]), .QN());
   DFF_X1 \values_reg[43][12]  (.D(values[12]), .CK(n_121_76), .Q(
      \values[43] [12]), .QN());
   DFF_X1 \values_reg[43][11]  (.D(values[11]), .CK(n_121_76), .Q(
      \values[43] [11]), .QN());
   DFF_X1 \values_reg[43][10]  (.D(values[10]), .CK(n_121_76), .Q(
      \values[43] [10]), .QN());
   DFF_X1 \values_reg[43][9]  (.D(values[9]), .CK(n_121_76), .Q(\values[43] [9]), 
      .QN());
   DFF_X1 \values_reg[43][8]  (.D(values[8]), .CK(n_121_76), .Q(\values[43] [8]), 
      .QN());
   DFF_X1 \values_reg[43][7]  (.D(values[7]), .CK(n_121_76), .Q(\values[43] [7]), 
      .QN());
   DFF_X1 \values_reg[43][6]  (.D(values[6]), .CK(n_121_76), .Q(\values[43] [6]), 
      .QN());
   DFF_X1 \values_reg[43][5]  (.D(values[5]), .CK(n_121_76), .Q(\values[43] [5]), 
      .QN());
   DFF_X1 \values_reg[43][4]  (.D(values[4]), .CK(n_121_76), .Q(\values[43] [4]), 
      .QN());
   DFF_X1 \values_reg[43][3]  (.D(values[3]), .CK(n_121_76), .Q(\values[43] [3]), 
      .QN());
   DFF_X1 \values_reg[43][2]  (.D(values[2]), .CK(n_121_76), .Q(\values[43] [2]), 
      .QN());
   DFF_X1 \values_reg[43][1]  (.D(values[1]), .CK(n_121_76), .Q(\values[43] [1]), 
      .QN());
   DFF_X1 \values_reg[43][0]  (.D(values[0]), .CK(n_121_76), .Q(\values[43] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[42]_reg  (.CK(clk), .E(n_42), .SE(1'b0), 
      .GCK(n_121_77));
   DFF_X1 \values_reg[42][15]  (.D(values[15]), .CK(n_121_77), .Q(
      \values[42] [15]), .QN());
   DFF_X1 \values_reg[42][14]  (.D(values[14]), .CK(n_121_77), .Q(
      \values[42] [14]), .QN());
   DFF_X1 \values_reg[42][13]  (.D(values[13]), .CK(n_121_77), .Q(
      \values[42] [13]), .QN());
   DFF_X1 \values_reg[42][12]  (.D(values[12]), .CK(n_121_77), .Q(
      \values[42] [12]), .QN());
   DFF_X1 \values_reg[42][11]  (.D(values[11]), .CK(n_121_77), .Q(
      \values[42] [11]), .QN());
   DFF_X1 \values_reg[42][10]  (.D(values[10]), .CK(n_121_77), .Q(
      \values[42] [10]), .QN());
   DFF_X1 \values_reg[42][9]  (.D(values[9]), .CK(n_121_77), .Q(\values[42] [9]), 
      .QN());
   DFF_X1 \values_reg[42][8]  (.D(values[8]), .CK(n_121_77), .Q(\values[42] [8]), 
      .QN());
   DFF_X1 \values_reg[42][7]  (.D(values[7]), .CK(n_121_77), .Q(\values[42] [7]), 
      .QN());
   DFF_X1 \values_reg[42][6]  (.D(values[6]), .CK(n_121_77), .Q(\values[42] [6]), 
      .QN());
   DFF_X1 \values_reg[42][5]  (.D(values[5]), .CK(n_121_77), .Q(\values[42] [5]), 
      .QN());
   DFF_X1 \values_reg[42][4]  (.D(values[4]), .CK(n_121_77), .Q(\values[42] [4]), 
      .QN());
   DFF_X1 \values_reg[42][3]  (.D(values[3]), .CK(n_121_77), .Q(\values[42] [3]), 
      .QN());
   DFF_X1 \values_reg[42][2]  (.D(values[2]), .CK(n_121_77), .Q(\values[42] [2]), 
      .QN());
   DFF_X1 \values_reg[42][1]  (.D(values[1]), .CK(n_121_77), .Q(\values[42] [1]), 
      .QN());
   DFF_X1 \values_reg[42][0]  (.D(values[0]), .CK(n_121_77), .Q(\values[42] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[41]_reg  (.CK(clk), .E(n_41), .SE(1'b0), 
      .GCK(n_121_78));
   DFF_X1 \values_reg[41][15]  (.D(values[15]), .CK(n_121_78), .Q(
      \values[41] [15]), .QN());
   DFF_X1 \values_reg[41][14]  (.D(values[14]), .CK(n_121_78), .Q(
      \values[41] [14]), .QN());
   DFF_X1 \values_reg[41][13]  (.D(values[13]), .CK(n_121_78), .Q(
      \values[41] [13]), .QN());
   DFF_X1 \values_reg[41][12]  (.D(values[12]), .CK(n_121_78), .Q(
      \values[41] [12]), .QN());
   DFF_X1 \values_reg[41][11]  (.D(values[11]), .CK(n_121_78), .Q(
      \values[41] [11]), .QN());
   DFF_X1 \values_reg[41][10]  (.D(values[10]), .CK(n_121_78), .Q(
      \values[41] [10]), .QN());
   DFF_X1 \values_reg[41][9]  (.D(values[9]), .CK(n_121_78), .Q(\values[41] [9]), 
      .QN());
   DFF_X1 \values_reg[41][8]  (.D(values[8]), .CK(n_121_78), .Q(\values[41] [8]), 
      .QN());
   DFF_X1 \values_reg[41][7]  (.D(values[7]), .CK(n_121_78), .Q(\values[41] [7]), 
      .QN());
   DFF_X1 \values_reg[41][6]  (.D(values[6]), .CK(n_121_78), .Q(\values[41] [6]), 
      .QN());
   DFF_X1 \values_reg[41][5]  (.D(values[5]), .CK(n_121_78), .Q(\values[41] [5]), 
      .QN());
   DFF_X1 \values_reg[41][4]  (.D(values[4]), .CK(n_121_78), .Q(\values[41] [4]), 
      .QN());
   DFF_X1 \values_reg[41][3]  (.D(values[3]), .CK(n_121_78), .Q(\values[41] [3]), 
      .QN());
   DFF_X1 \values_reg[41][2]  (.D(values[2]), .CK(n_121_78), .Q(\values[41] [2]), 
      .QN());
   DFF_X1 \values_reg[41][1]  (.D(values[1]), .CK(n_121_78), .Q(\values[41] [1]), 
      .QN());
   DFF_X1 \values_reg[41][0]  (.D(values[0]), .CK(n_121_78), .Q(\values[41] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[40]_reg  (.CK(clk), .E(n_40), .SE(1'b0), 
      .GCK(n_121_79));
   DFF_X1 \values_reg[40][15]  (.D(values[15]), .CK(n_121_79), .Q(
      \values[40] [15]), .QN());
   DFF_X1 \values_reg[40][14]  (.D(values[14]), .CK(n_121_79), .Q(
      \values[40] [14]), .QN());
   DFF_X1 \values_reg[40][13]  (.D(values[13]), .CK(n_121_79), .Q(
      \values[40] [13]), .QN());
   DFF_X1 \values_reg[40][12]  (.D(values[12]), .CK(n_121_79), .Q(
      \values[40] [12]), .QN());
   DFF_X1 \values_reg[40][11]  (.D(values[11]), .CK(n_121_79), .Q(
      \values[40] [11]), .QN());
   DFF_X1 \values_reg[40][10]  (.D(values[10]), .CK(n_121_79), .Q(
      \values[40] [10]), .QN());
   DFF_X1 \values_reg[40][9]  (.D(values[9]), .CK(n_121_79), .Q(\values[40] [9]), 
      .QN());
   DFF_X1 \values_reg[40][8]  (.D(values[8]), .CK(n_121_79), .Q(\values[40] [8]), 
      .QN());
   DFF_X1 \values_reg[40][7]  (.D(values[7]), .CK(n_121_79), .Q(\values[40] [7]), 
      .QN());
   DFF_X1 \values_reg[40][6]  (.D(values[6]), .CK(n_121_79), .Q(\values[40] [6]), 
      .QN());
   DFF_X1 \values_reg[40][5]  (.D(values[5]), .CK(n_121_79), .Q(\values[40] [5]), 
      .QN());
   DFF_X1 \values_reg[40][4]  (.D(values[4]), .CK(n_121_79), .Q(\values[40] [4]), 
      .QN());
   DFF_X1 \values_reg[40][3]  (.D(values[3]), .CK(n_121_79), .Q(\values[40] [3]), 
      .QN());
   DFF_X1 \values_reg[40][2]  (.D(values[2]), .CK(n_121_79), .Q(\values[40] [2]), 
      .QN());
   DFF_X1 \values_reg[40][1]  (.D(values[1]), .CK(n_121_79), .Q(\values[40] [1]), 
      .QN());
   DFF_X1 \values_reg[40][0]  (.D(values[0]), .CK(n_121_79), .Q(\values[40] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[39]_reg  (.CK(clk), .E(n_39), .SE(1'b0), 
      .GCK(n_121_80));
   DFF_X1 \values_reg[39][15]  (.D(values[15]), .CK(n_121_80), .Q(
      \values[39] [15]), .QN());
   DFF_X1 \values_reg[39][14]  (.D(values[14]), .CK(n_121_80), .Q(
      \values[39] [14]), .QN());
   DFF_X1 \values_reg[39][13]  (.D(values[13]), .CK(n_121_80), .Q(
      \values[39] [13]), .QN());
   DFF_X1 \values_reg[39][12]  (.D(values[12]), .CK(n_121_80), .Q(
      \values[39] [12]), .QN());
   DFF_X1 \values_reg[39][11]  (.D(values[11]), .CK(n_121_80), .Q(
      \values[39] [11]), .QN());
   DFF_X1 \values_reg[39][10]  (.D(values[10]), .CK(n_121_80), .Q(
      \values[39] [10]), .QN());
   DFF_X1 \values_reg[39][9]  (.D(values[9]), .CK(n_121_80), .Q(\values[39] [9]), 
      .QN());
   DFF_X1 \values_reg[39][8]  (.D(values[8]), .CK(n_121_80), .Q(\values[39] [8]), 
      .QN());
   DFF_X1 \values_reg[39][7]  (.D(values[7]), .CK(n_121_80), .Q(\values[39] [7]), 
      .QN());
   DFF_X1 \values_reg[39][6]  (.D(values[6]), .CK(n_121_80), .Q(\values[39] [6]), 
      .QN());
   DFF_X1 \values_reg[39][5]  (.D(values[5]), .CK(n_121_80), .Q(\values[39] [5]), 
      .QN());
   DFF_X1 \values_reg[39][4]  (.D(values[4]), .CK(n_121_80), .Q(\values[39] [4]), 
      .QN());
   DFF_X1 \values_reg[39][3]  (.D(values[3]), .CK(n_121_80), .Q(\values[39] [3]), 
      .QN());
   DFF_X1 \values_reg[39][2]  (.D(values[2]), .CK(n_121_80), .Q(\values[39] [2]), 
      .QN());
   DFF_X1 \values_reg[39][1]  (.D(values[1]), .CK(n_121_80), .Q(\values[39] [1]), 
      .QN());
   DFF_X1 \values_reg[39][0]  (.D(values[0]), .CK(n_121_80), .Q(\values[39] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[38]_reg  (.CK(clk), .E(n_38), .SE(1'b0), 
      .GCK(n_121_81));
   DFF_X1 \values_reg[38][15]  (.D(values[15]), .CK(n_121_81), .Q(
      \values[38] [15]), .QN());
   DFF_X1 \values_reg[38][14]  (.D(values[14]), .CK(n_121_81), .Q(
      \values[38] [14]), .QN());
   DFF_X1 \values_reg[38][13]  (.D(values[13]), .CK(n_121_81), .Q(
      \values[38] [13]), .QN());
   DFF_X1 \values_reg[38][12]  (.D(values[12]), .CK(n_121_81), .Q(
      \values[38] [12]), .QN());
   DFF_X1 \values_reg[38][11]  (.D(values[11]), .CK(n_121_81), .Q(
      \values[38] [11]), .QN());
   DFF_X1 \values_reg[38][10]  (.D(values[10]), .CK(n_121_81), .Q(
      \values[38] [10]), .QN());
   DFF_X1 \values_reg[38][9]  (.D(values[9]), .CK(n_121_81), .Q(\values[38] [9]), 
      .QN());
   DFF_X1 \values_reg[38][8]  (.D(values[8]), .CK(n_121_81), .Q(\values[38] [8]), 
      .QN());
   DFF_X1 \values_reg[38][7]  (.D(values[7]), .CK(n_121_81), .Q(\values[38] [7]), 
      .QN());
   DFF_X1 \values_reg[38][6]  (.D(values[6]), .CK(n_121_81), .Q(\values[38] [6]), 
      .QN());
   DFF_X1 \values_reg[38][5]  (.D(values[5]), .CK(n_121_81), .Q(\values[38] [5]), 
      .QN());
   DFF_X1 \values_reg[38][4]  (.D(values[4]), .CK(n_121_81), .Q(\values[38] [4]), 
      .QN());
   DFF_X1 \values_reg[38][3]  (.D(values[3]), .CK(n_121_81), .Q(\values[38] [3]), 
      .QN());
   DFF_X1 \values_reg[38][2]  (.D(values[2]), .CK(n_121_81), .Q(\values[38] [2]), 
      .QN());
   DFF_X1 \values_reg[38][1]  (.D(values[1]), .CK(n_121_81), .Q(\values[38] [1]), 
      .QN());
   DFF_X1 \values_reg[38][0]  (.D(values[0]), .CK(n_121_81), .Q(\values[38] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[37]_reg  (.CK(clk), .E(n_37), .SE(1'b0), 
      .GCK(n_121_82));
   DFF_X1 \values_reg[37][15]  (.D(values[15]), .CK(n_121_82), .Q(
      \values[37] [15]), .QN());
   DFF_X1 \values_reg[37][14]  (.D(values[14]), .CK(n_121_82), .Q(
      \values[37] [14]), .QN());
   DFF_X1 \values_reg[37][13]  (.D(values[13]), .CK(n_121_82), .Q(
      \values[37] [13]), .QN());
   DFF_X1 \values_reg[37][12]  (.D(values[12]), .CK(n_121_82), .Q(
      \values[37] [12]), .QN());
   DFF_X1 \values_reg[37][11]  (.D(values[11]), .CK(n_121_82), .Q(
      \values[37] [11]), .QN());
   DFF_X1 \values_reg[37][10]  (.D(values[10]), .CK(n_121_82), .Q(
      \values[37] [10]), .QN());
   DFF_X1 \values_reg[37][9]  (.D(values[9]), .CK(n_121_82), .Q(\values[37] [9]), 
      .QN());
   DFF_X1 \values_reg[37][8]  (.D(values[8]), .CK(n_121_82), .Q(\values[37] [8]), 
      .QN());
   DFF_X1 \values_reg[37][7]  (.D(values[7]), .CK(n_121_82), .Q(\values[37] [7]), 
      .QN());
   DFF_X1 \values_reg[37][6]  (.D(values[6]), .CK(n_121_82), .Q(\values[37] [6]), 
      .QN());
   DFF_X1 \values_reg[37][5]  (.D(values[5]), .CK(n_121_82), .Q(\values[37] [5]), 
      .QN());
   DFF_X1 \values_reg[37][4]  (.D(values[4]), .CK(n_121_82), .Q(\values[37] [4]), 
      .QN());
   DFF_X1 \values_reg[37][3]  (.D(values[3]), .CK(n_121_82), .Q(\values[37] [3]), 
      .QN());
   DFF_X1 \values_reg[37][2]  (.D(values[2]), .CK(n_121_82), .Q(\values[37] [2]), 
      .QN());
   DFF_X1 \values_reg[37][1]  (.D(values[1]), .CK(n_121_82), .Q(\values[37] [1]), 
      .QN());
   DFF_X1 \values_reg[37][0]  (.D(values[0]), .CK(n_121_82), .Q(\values[37] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[36]_reg  (.CK(clk), .E(n_36), .SE(1'b0), 
      .GCK(n_121_83));
   DFF_X1 \values_reg[36][15]  (.D(values[15]), .CK(n_121_83), .Q(
      \values[36] [15]), .QN());
   DFF_X1 \values_reg[36][14]  (.D(values[14]), .CK(n_121_83), .Q(
      \values[36] [14]), .QN());
   DFF_X1 \values_reg[36][13]  (.D(values[13]), .CK(n_121_83), .Q(
      \values[36] [13]), .QN());
   DFF_X1 \values_reg[36][12]  (.D(values[12]), .CK(n_121_83), .Q(
      \values[36] [12]), .QN());
   DFF_X1 \values_reg[36][11]  (.D(values[11]), .CK(n_121_83), .Q(
      \values[36] [11]), .QN());
   DFF_X1 \values_reg[36][10]  (.D(values[10]), .CK(n_121_83), .Q(
      \values[36] [10]), .QN());
   DFF_X1 \values_reg[36][9]  (.D(values[9]), .CK(n_121_83), .Q(\values[36] [9]), 
      .QN());
   DFF_X1 \values_reg[36][8]  (.D(values[8]), .CK(n_121_83), .Q(\values[36] [8]), 
      .QN());
   DFF_X1 \values_reg[36][7]  (.D(values[7]), .CK(n_121_83), .Q(\values[36] [7]), 
      .QN());
   DFF_X1 \values_reg[36][6]  (.D(values[6]), .CK(n_121_83), .Q(\values[36] [6]), 
      .QN());
   DFF_X1 \values_reg[36][5]  (.D(values[5]), .CK(n_121_83), .Q(\values[36] [5]), 
      .QN());
   DFF_X1 \values_reg[36][4]  (.D(values[4]), .CK(n_121_83), .Q(\values[36] [4]), 
      .QN());
   DFF_X1 \values_reg[36][3]  (.D(values[3]), .CK(n_121_83), .Q(\values[36] [3]), 
      .QN());
   DFF_X1 \values_reg[36][2]  (.D(values[2]), .CK(n_121_83), .Q(\values[36] [2]), 
      .QN());
   DFF_X1 \values_reg[36][1]  (.D(values[1]), .CK(n_121_83), .Q(\values[36] [1]), 
      .QN());
   DFF_X1 \values_reg[36][0]  (.D(values[0]), .CK(n_121_83), .Q(\values[36] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[35]_reg  (.CK(clk), .E(n_35), .SE(1'b0), 
      .GCK(n_121_84));
   DFF_X1 \values_reg[35][15]  (.D(values[15]), .CK(n_121_84), .Q(
      \values[35] [15]), .QN());
   DFF_X1 \values_reg[35][14]  (.D(values[14]), .CK(n_121_84), .Q(
      \values[35] [14]), .QN());
   DFF_X1 \values_reg[35][13]  (.D(values[13]), .CK(n_121_84), .Q(
      \values[35] [13]), .QN());
   DFF_X1 \values_reg[35][12]  (.D(values[12]), .CK(n_121_84), .Q(
      \values[35] [12]), .QN());
   DFF_X1 \values_reg[35][11]  (.D(values[11]), .CK(n_121_84), .Q(
      \values[35] [11]), .QN());
   DFF_X1 \values_reg[35][10]  (.D(values[10]), .CK(n_121_84), .Q(
      \values[35] [10]), .QN());
   DFF_X1 \values_reg[35][9]  (.D(values[9]), .CK(n_121_84), .Q(\values[35] [9]), 
      .QN());
   DFF_X1 \values_reg[35][8]  (.D(values[8]), .CK(n_121_84), .Q(\values[35] [8]), 
      .QN());
   DFF_X1 \values_reg[35][7]  (.D(values[7]), .CK(n_121_84), .Q(\values[35] [7]), 
      .QN());
   DFF_X1 \values_reg[35][6]  (.D(values[6]), .CK(n_121_84), .Q(\values[35] [6]), 
      .QN());
   DFF_X1 \values_reg[35][5]  (.D(values[5]), .CK(n_121_84), .Q(\values[35] [5]), 
      .QN());
   DFF_X1 \values_reg[35][4]  (.D(values[4]), .CK(n_121_84), .Q(\values[35] [4]), 
      .QN());
   DFF_X1 \values_reg[35][3]  (.D(values[3]), .CK(n_121_84), .Q(\values[35] [3]), 
      .QN());
   DFF_X1 \values_reg[35][2]  (.D(values[2]), .CK(n_121_84), .Q(\values[35] [2]), 
      .QN());
   DFF_X1 \values_reg[35][1]  (.D(values[1]), .CK(n_121_84), .Q(\values[35] [1]), 
      .QN());
   DFF_X1 \values_reg[35][0]  (.D(values[0]), .CK(n_121_84), .Q(\values[35] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[34]_reg  (.CK(clk), .E(n_34), .SE(1'b0), 
      .GCK(n_121_85));
   DFF_X1 \values_reg[34][15]  (.D(values[15]), .CK(n_121_85), .Q(
      \values[34] [15]), .QN());
   DFF_X1 \values_reg[34][14]  (.D(values[14]), .CK(n_121_85), .Q(
      \values[34] [14]), .QN());
   DFF_X1 \values_reg[34][13]  (.D(values[13]), .CK(n_121_85), .Q(
      \values[34] [13]), .QN());
   DFF_X1 \values_reg[34][12]  (.D(values[12]), .CK(n_121_85), .Q(
      \values[34] [12]), .QN());
   DFF_X1 \values_reg[34][11]  (.D(values[11]), .CK(n_121_85), .Q(
      \values[34] [11]), .QN());
   DFF_X1 \values_reg[34][10]  (.D(values[10]), .CK(n_121_85), .Q(
      \values[34] [10]), .QN());
   DFF_X1 \values_reg[34][9]  (.D(values[9]), .CK(n_121_85), .Q(\values[34] [9]), 
      .QN());
   DFF_X1 \values_reg[34][8]  (.D(values[8]), .CK(n_121_85), .Q(\values[34] [8]), 
      .QN());
   DFF_X1 \values_reg[34][7]  (.D(values[7]), .CK(n_121_85), .Q(\values[34] [7]), 
      .QN());
   DFF_X1 \values_reg[34][6]  (.D(values[6]), .CK(n_121_85), .Q(\values[34] [6]), 
      .QN());
   DFF_X1 \values_reg[34][5]  (.D(values[5]), .CK(n_121_85), .Q(\values[34] [5]), 
      .QN());
   DFF_X1 \values_reg[34][4]  (.D(values[4]), .CK(n_121_85), .Q(\values[34] [4]), 
      .QN());
   DFF_X1 \values_reg[34][3]  (.D(values[3]), .CK(n_121_85), .Q(\values[34] [3]), 
      .QN());
   DFF_X1 \values_reg[34][2]  (.D(values[2]), .CK(n_121_85), .Q(\values[34] [2]), 
      .QN());
   DFF_X1 \values_reg[34][1]  (.D(values[1]), .CK(n_121_85), .Q(\values[34] [1]), 
      .QN());
   DFF_X1 \values_reg[34][0]  (.D(values[0]), .CK(n_121_85), .Q(\values[34] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[33]_reg  (.CK(clk), .E(n_33), .SE(1'b0), 
      .GCK(n_121_86));
   DFF_X1 \values_reg[33][15]  (.D(values[15]), .CK(n_121_86), .Q(
      \values[33] [15]), .QN());
   DFF_X1 \values_reg[33][14]  (.D(values[14]), .CK(n_121_86), .Q(
      \values[33] [14]), .QN());
   DFF_X1 \values_reg[33][13]  (.D(values[13]), .CK(n_121_86), .Q(
      \values[33] [13]), .QN());
   DFF_X1 \values_reg[33][12]  (.D(values[12]), .CK(n_121_86), .Q(
      \values[33] [12]), .QN());
   DFF_X1 \values_reg[33][11]  (.D(values[11]), .CK(n_121_86), .Q(
      \values[33] [11]), .QN());
   DFF_X1 \values_reg[33][10]  (.D(values[10]), .CK(n_121_86), .Q(
      \values[33] [10]), .QN());
   DFF_X1 \values_reg[33][9]  (.D(values[9]), .CK(n_121_86), .Q(\values[33] [9]), 
      .QN());
   DFF_X1 \values_reg[33][8]  (.D(values[8]), .CK(n_121_86), .Q(\values[33] [8]), 
      .QN());
   DFF_X1 \values_reg[33][7]  (.D(values[7]), .CK(n_121_86), .Q(\values[33] [7]), 
      .QN());
   DFF_X1 \values_reg[33][6]  (.D(values[6]), .CK(n_121_86), .Q(\values[33] [6]), 
      .QN());
   DFF_X1 \values_reg[33][5]  (.D(values[5]), .CK(n_121_86), .Q(\values[33] [5]), 
      .QN());
   DFF_X1 \values_reg[33][4]  (.D(values[4]), .CK(n_121_86), .Q(\values[33] [4]), 
      .QN());
   DFF_X1 \values_reg[33][3]  (.D(values[3]), .CK(n_121_86), .Q(\values[33] [3]), 
      .QN());
   DFF_X1 \values_reg[33][2]  (.D(values[2]), .CK(n_121_86), .Q(\values[33] [2]), 
      .QN());
   DFF_X1 \values_reg[33][1]  (.D(values[1]), .CK(n_121_86), .Q(\values[33] [1]), 
      .QN());
   DFF_X1 \values_reg[33][0]  (.D(values[0]), .CK(n_121_86), .Q(\values[33] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[32]_reg  (.CK(clk), .E(n_32), .SE(1'b0), 
      .GCK(n_121_87));
   DFF_X1 \values_reg[32][15]  (.D(values[15]), .CK(n_121_87), .Q(
      \values[32] [15]), .QN());
   DFF_X1 \values_reg[32][14]  (.D(values[14]), .CK(n_121_87), .Q(
      \values[32] [14]), .QN());
   DFF_X1 \values_reg[32][13]  (.D(values[13]), .CK(n_121_87), .Q(
      \values[32] [13]), .QN());
   DFF_X1 \values_reg[32][12]  (.D(values[12]), .CK(n_121_87), .Q(
      \values[32] [12]), .QN());
   DFF_X1 \values_reg[32][11]  (.D(values[11]), .CK(n_121_87), .Q(
      \values[32] [11]), .QN());
   DFF_X1 \values_reg[32][10]  (.D(values[10]), .CK(n_121_87), .Q(
      \values[32] [10]), .QN());
   DFF_X1 \values_reg[32][9]  (.D(values[9]), .CK(n_121_87), .Q(\values[32] [9]), 
      .QN());
   DFF_X1 \values_reg[32][8]  (.D(values[8]), .CK(n_121_87), .Q(\values[32] [8]), 
      .QN());
   DFF_X1 \values_reg[32][7]  (.D(values[7]), .CK(n_121_87), .Q(\values[32] [7]), 
      .QN());
   DFF_X1 \values_reg[32][6]  (.D(values[6]), .CK(n_121_87), .Q(\values[32] [6]), 
      .QN());
   DFF_X1 \values_reg[32][5]  (.D(values[5]), .CK(n_121_87), .Q(\values[32] [5]), 
      .QN());
   DFF_X1 \values_reg[32][4]  (.D(values[4]), .CK(n_121_87), .Q(\values[32] [4]), 
      .QN());
   DFF_X1 \values_reg[32][3]  (.D(values[3]), .CK(n_121_87), .Q(\values[32] [3]), 
      .QN());
   DFF_X1 \values_reg[32][2]  (.D(values[2]), .CK(n_121_87), .Q(\values[32] [2]), 
      .QN());
   DFF_X1 \values_reg[32][1]  (.D(values[1]), .CK(n_121_87), .Q(\values[32] [1]), 
      .QN());
   DFF_X1 \values_reg[32][0]  (.D(values[0]), .CK(n_121_87), .Q(\values[32] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[31]_reg  (.CK(clk), .E(n_31), .SE(1'b0), 
      .GCK(n_121_88));
   DFF_X1 \values_reg[31][15]  (.D(values[15]), .CK(n_121_88), .Q(
      \values[31] [15]), .QN());
   DFF_X1 \values_reg[31][14]  (.D(values[14]), .CK(n_121_88), .Q(
      \values[31] [14]), .QN());
   DFF_X1 \values_reg[31][13]  (.D(values[13]), .CK(n_121_88), .Q(
      \values[31] [13]), .QN());
   DFF_X1 \values_reg[31][12]  (.D(values[12]), .CK(n_121_88), .Q(
      \values[31] [12]), .QN());
   DFF_X1 \values_reg[31][11]  (.D(values[11]), .CK(n_121_88), .Q(
      \values[31] [11]), .QN());
   DFF_X1 \values_reg[31][10]  (.D(values[10]), .CK(n_121_88), .Q(
      \values[31] [10]), .QN());
   DFF_X1 \values_reg[31][9]  (.D(values[9]), .CK(n_121_88), .Q(\values[31] [9]), 
      .QN());
   DFF_X1 \values_reg[31][8]  (.D(values[8]), .CK(n_121_88), .Q(\values[31] [8]), 
      .QN());
   DFF_X1 \values_reg[31][7]  (.D(values[7]), .CK(n_121_88), .Q(\values[31] [7]), 
      .QN());
   DFF_X1 \values_reg[31][6]  (.D(values[6]), .CK(n_121_88), .Q(\values[31] [6]), 
      .QN());
   DFF_X1 \values_reg[31][5]  (.D(values[5]), .CK(n_121_88), .Q(\values[31] [5]), 
      .QN());
   DFF_X1 \values_reg[31][4]  (.D(values[4]), .CK(n_121_88), .Q(\values[31] [4]), 
      .QN());
   DFF_X1 \values_reg[31][3]  (.D(values[3]), .CK(n_121_88), .Q(\values[31] [3]), 
      .QN());
   DFF_X1 \values_reg[31][2]  (.D(values[2]), .CK(n_121_88), .Q(\values[31] [2]), 
      .QN());
   DFF_X1 \values_reg[31][1]  (.D(values[1]), .CK(n_121_88), .Q(\values[31] [1]), 
      .QN());
   DFF_X1 \values_reg[31][0]  (.D(values[0]), .CK(n_121_88), .Q(\values[31] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[30]_reg  (.CK(clk), .E(n_30), .SE(1'b0), 
      .GCK(n_121_89));
   DFF_X1 \values_reg[30][15]  (.D(values[15]), .CK(n_121_89), .Q(
      \values[30] [15]), .QN());
   DFF_X1 \values_reg[30][14]  (.D(values[14]), .CK(n_121_89), .Q(
      \values[30] [14]), .QN());
   DFF_X1 \values_reg[30][13]  (.D(values[13]), .CK(n_121_89), .Q(
      \values[30] [13]), .QN());
   DFF_X1 \values_reg[30][12]  (.D(values[12]), .CK(n_121_89), .Q(
      \values[30] [12]), .QN());
   DFF_X1 \values_reg[30][11]  (.D(values[11]), .CK(n_121_89), .Q(
      \values[30] [11]), .QN());
   DFF_X1 \values_reg[30][10]  (.D(values[10]), .CK(n_121_89), .Q(
      \values[30] [10]), .QN());
   DFF_X1 \values_reg[30][9]  (.D(values[9]), .CK(n_121_89), .Q(\values[30] [9]), 
      .QN());
   DFF_X1 \values_reg[30][8]  (.D(values[8]), .CK(n_121_89), .Q(\values[30] [8]), 
      .QN());
   DFF_X1 \values_reg[30][7]  (.D(values[7]), .CK(n_121_89), .Q(\values[30] [7]), 
      .QN());
   DFF_X1 \values_reg[30][6]  (.D(values[6]), .CK(n_121_89), .Q(\values[30] [6]), 
      .QN());
   DFF_X1 \values_reg[30][5]  (.D(values[5]), .CK(n_121_89), .Q(\values[30] [5]), 
      .QN());
   DFF_X1 \values_reg[30][4]  (.D(values[4]), .CK(n_121_89), .Q(\values[30] [4]), 
      .QN());
   DFF_X1 \values_reg[30][3]  (.D(values[3]), .CK(n_121_89), .Q(\values[30] [3]), 
      .QN());
   DFF_X1 \values_reg[30][2]  (.D(values[2]), .CK(n_121_89), .Q(\values[30] [2]), 
      .QN());
   DFF_X1 \values_reg[30][1]  (.D(values[1]), .CK(n_121_89), .Q(\values[30] [1]), 
      .QN());
   DFF_X1 \values_reg[30][0]  (.D(values[0]), .CK(n_121_89), .Q(\values[30] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[29]_reg  (.CK(clk), .E(n_29), .SE(1'b0), 
      .GCK(n_121_90));
   DFF_X1 \values_reg[29][15]  (.D(values[15]), .CK(n_121_90), .Q(
      \values[29] [15]), .QN());
   DFF_X1 \values_reg[29][14]  (.D(values[14]), .CK(n_121_90), .Q(
      \values[29] [14]), .QN());
   DFF_X1 \values_reg[29][13]  (.D(values[13]), .CK(n_121_90), .Q(
      \values[29] [13]), .QN());
   DFF_X1 \values_reg[29][12]  (.D(values[12]), .CK(n_121_90), .Q(
      \values[29] [12]), .QN());
   DFF_X1 \values_reg[29][11]  (.D(values[11]), .CK(n_121_90), .Q(
      \values[29] [11]), .QN());
   DFF_X1 \values_reg[29][10]  (.D(values[10]), .CK(n_121_90), .Q(
      \values[29] [10]), .QN());
   DFF_X1 \values_reg[29][9]  (.D(values[9]), .CK(n_121_90), .Q(\values[29] [9]), 
      .QN());
   DFF_X1 \values_reg[29][8]  (.D(values[8]), .CK(n_121_90), .Q(\values[29] [8]), 
      .QN());
   DFF_X1 \values_reg[29][7]  (.D(values[7]), .CK(n_121_90), .Q(\values[29] [7]), 
      .QN());
   DFF_X1 \values_reg[29][6]  (.D(values[6]), .CK(n_121_90), .Q(\values[29] [6]), 
      .QN());
   DFF_X1 \values_reg[29][5]  (.D(values[5]), .CK(n_121_90), .Q(\values[29] [5]), 
      .QN());
   DFF_X1 \values_reg[29][4]  (.D(values[4]), .CK(n_121_90), .Q(\values[29] [4]), 
      .QN());
   DFF_X1 \values_reg[29][3]  (.D(values[3]), .CK(n_121_90), .Q(\values[29] [3]), 
      .QN());
   DFF_X1 \values_reg[29][2]  (.D(values[2]), .CK(n_121_90), .Q(\values[29] [2]), 
      .QN());
   DFF_X1 \values_reg[29][1]  (.D(values[1]), .CK(n_121_90), .Q(\values[29] [1]), 
      .QN());
   DFF_X1 \values_reg[29][0]  (.D(values[0]), .CK(n_121_90), .Q(\values[29] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[28]_reg  (.CK(clk), .E(n_28), .SE(1'b0), 
      .GCK(n_121_91));
   DFF_X1 \values_reg[28][15]  (.D(values[15]), .CK(n_121_91), .Q(
      \values[28] [15]), .QN());
   DFF_X1 \values_reg[28][14]  (.D(values[14]), .CK(n_121_91), .Q(
      \values[28] [14]), .QN());
   DFF_X1 \values_reg[28][13]  (.D(values[13]), .CK(n_121_91), .Q(
      \values[28] [13]), .QN());
   DFF_X1 \values_reg[28][12]  (.D(values[12]), .CK(n_121_91), .Q(
      \values[28] [12]), .QN());
   DFF_X1 \values_reg[28][11]  (.D(values[11]), .CK(n_121_91), .Q(
      \values[28] [11]), .QN());
   DFF_X1 \values_reg[28][10]  (.D(values[10]), .CK(n_121_91), .Q(
      \values[28] [10]), .QN());
   DFF_X1 \values_reg[28][9]  (.D(values[9]), .CK(n_121_91), .Q(\values[28] [9]), 
      .QN());
   DFF_X1 \values_reg[28][8]  (.D(values[8]), .CK(n_121_91), .Q(\values[28] [8]), 
      .QN());
   DFF_X1 \values_reg[28][7]  (.D(values[7]), .CK(n_121_91), .Q(\values[28] [7]), 
      .QN());
   DFF_X1 \values_reg[28][6]  (.D(values[6]), .CK(n_121_91), .Q(\values[28] [6]), 
      .QN());
   DFF_X1 \values_reg[28][5]  (.D(values[5]), .CK(n_121_91), .Q(\values[28] [5]), 
      .QN());
   DFF_X1 \values_reg[28][4]  (.D(values[4]), .CK(n_121_91), .Q(\values[28] [4]), 
      .QN());
   DFF_X1 \values_reg[28][3]  (.D(values[3]), .CK(n_121_91), .Q(\values[28] [3]), 
      .QN());
   DFF_X1 \values_reg[28][2]  (.D(values[2]), .CK(n_121_91), .Q(\values[28] [2]), 
      .QN());
   DFF_X1 \values_reg[28][1]  (.D(values[1]), .CK(n_121_91), .Q(\values[28] [1]), 
      .QN());
   DFF_X1 \values_reg[28][0]  (.D(values[0]), .CK(n_121_91), .Q(\values[28] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[27]_reg  (.CK(clk), .E(n_27), .SE(1'b0), 
      .GCK(n_121_92));
   DFF_X1 \values_reg[27][15]  (.D(values[15]), .CK(n_121_92), .Q(
      \values[27] [15]), .QN());
   DFF_X1 \values_reg[27][14]  (.D(values[14]), .CK(n_121_92), .Q(
      \values[27] [14]), .QN());
   DFF_X1 \values_reg[27][13]  (.D(values[13]), .CK(n_121_92), .Q(
      \values[27] [13]), .QN());
   DFF_X1 \values_reg[27][12]  (.D(values[12]), .CK(n_121_92), .Q(
      \values[27] [12]), .QN());
   DFF_X1 \values_reg[27][11]  (.D(values[11]), .CK(n_121_92), .Q(
      \values[27] [11]), .QN());
   DFF_X1 \values_reg[27][10]  (.D(values[10]), .CK(n_121_92), .Q(
      \values[27] [10]), .QN());
   DFF_X1 \values_reg[27][9]  (.D(values[9]), .CK(n_121_92), .Q(\values[27] [9]), 
      .QN());
   DFF_X1 \values_reg[27][8]  (.D(values[8]), .CK(n_121_92), .Q(\values[27] [8]), 
      .QN());
   DFF_X1 \values_reg[27][7]  (.D(values[7]), .CK(n_121_92), .Q(\values[27] [7]), 
      .QN());
   DFF_X1 \values_reg[27][6]  (.D(values[6]), .CK(n_121_92), .Q(\values[27] [6]), 
      .QN());
   DFF_X1 \values_reg[27][5]  (.D(values[5]), .CK(n_121_92), .Q(\values[27] [5]), 
      .QN());
   DFF_X1 \values_reg[27][4]  (.D(values[4]), .CK(n_121_92), .Q(\values[27] [4]), 
      .QN());
   DFF_X1 \values_reg[27][3]  (.D(values[3]), .CK(n_121_92), .Q(\values[27] [3]), 
      .QN());
   DFF_X1 \values_reg[27][2]  (.D(values[2]), .CK(n_121_92), .Q(\values[27] [2]), 
      .QN());
   DFF_X1 \values_reg[27][1]  (.D(values[1]), .CK(n_121_92), .Q(\values[27] [1]), 
      .QN());
   DFF_X1 \values_reg[27][0]  (.D(values[0]), .CK(n_121_92), .Q(\values[27] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[26]_reg  (.CK(clk), .E(n_26), .SE(1'b0), 
      .GCK(n_121_93));
   DFF_X1 \values_reg[26][15]  (.D(values[15]), .CK(n_121_93), .Q(
      \values[26] [15]), .QN());
   DFF_X1 \values_reg[26][14]  (.D(values[14]), .CK(n_121_93), .Q(
      \values[26] [14]), .QN());
   DFF_X1 \values_reg[26][13]  (.D(values[13]), .CK(n_121_93), .Q(
      \values[26] [13]), .QN());
   DFF_X1 \values_reg[26][12]  (.D(values[12]), .CK(n_121_93), .Q(
      \values[26] [12]), .QN());
   DFF_X1 \values_reg[26][11]  (.D(values[11]), .CK(n_121_93), .Q(
      \values[26] [11]), .QN());
   DFF_X1 \values_reg[26][10]  (.D(values[10]), .CK(n_121_93), .Q(
      \values[26] [10]), .QN());
   DFF_X1 \values_reg[26][9]  (.D(values[9]), .CK(n_121_93), .Q(\values[26] [9]), 
      .QN());
   DFF_X1 \values_reg[26][8]  (.D(values[8]), .CK(n_121_93), .Q(\values[26] [8]), 
      .QN());
   DFF_X1 \values_reg[26][7]  (.D(values[7]), .CK(n_121_93), .Q(\values[26] [7]), 
      .QN());
   DFF_X1 \values_reg[26][6]  (.D(values[6]), .CK(n_121_93), .Q(\values[26] [6]), 
      .QN());
   DFF_X1 \values_reg[26][5]  (.D(values[5]), .CK(n_121_93), .Q(\values[26] [5]), 
      .QN());
   DFF_X1 \values_reg[26][4]  (.D(values[4]), .CK(n_121_93), .Q(\values[26] [4]), 
      .QN());
   DFF_X1 \values_reg[26][3]  (.D(values[3]), .CK(n_121_93), .Q(\values[26] [3]), 
      .QN());
   DFF_X1 \values_reg[26][2]  (.D(values[2]), .CK(n_121_93), .Q(\values[26] [2]), 
      .QN());
   DFF_X1 \values_reg[26][1]  (.D(values[1]), .CK(n_121_93), .Q(\values[26] [1]), 
      .QN());
   DFF_X1 \values_reg[26][0]  (.D(values[0]), .CK(n_121_93), .Q(\values[26] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[97]_reg  (.CK(clk), .E(n_97), .SE(1'b0), 
      .GCK(n_122_0));
   DFF_X1 \values_reg[97][15]  (.D(values[15]), .CK(n_122_0), .Q(
      \values[97] [15]), .QN());
   DFF_X1 \values_reg[97][14]  (.D(values[14]), .CK(n_122_0), .Q(
      \values[97] [14]), .QN());
   DFF_X1 \values_reg[97][13]  (.D(values[13]), .CK(n_122_0), .Q(
      \values[97] [13]), .QN());
   DFF_X1 \values_reg[97][12]  (.D(values[12]), .CK(n_122_0), .Q(
      \values[97] [12]), .QN());
   DFF_X1 \values_reg[97][11]  (.D(values[11]), .CK(n_122_0), .Q(
      \values[97] [11]), .QN());
   DFF_X1 \values_reg[97][10]  (.D(values[10]), .CK(n_122_0), .Q(
      \values[97] [10]), .QN());
   DFF_X1 \values_reg[97][9]  (.D(values[9]), .CK(n_122_0), .Q(\values[97] [9]), 
      .QN());
   DFF_X1 \values_reg[97][8]  (.D(values[8]), .CK(n_122_0), .Q(\values[97] [8]), 
      .QN());
   DFF_X1 \values_reg[97][7]  (.D(values[7]), .CK(n_122_0), .Q(\values[97] [7]), 
      .QN());
   DFF_X1 \values_reg[97][6]  (.D(values[6]), .CK(n_122_0), .Q(\values[97] [6]), 
      .QN());
   DFF_X1 \values_reg[97][5]  (.D(values[5]), .CK(n_122_0), .Q(\values[97] [5]), 
      .QN());
   DFF_X1 \values_reg[97][4]  (.D(values[4]), .CK(n_122_0), .Q(\values[97] [4]), 
      .QN());
   DFF_X1 \values_reg[97][3]  (.D(values[3]), .CK(n_122_0), .Q(\values[97] [3]), 
      .QN());
   DFF_X1 \values_reg[97][2]  (.D(values[2]), .CK(n_122_0), .Q(\values[97] [2]), 
      .QN());
   DFF_X1 \values_reg[97][1]  (.D(values[1]), .CK(n_122_0), .Q(\values[97] [1]), 
      .QN());
   DFF_X1 \values_reg[97][0]  (.D(values[0]), .CK(n_122_0), .Q(\values[97] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[98]_reg  (.CK(clk), .E(n_98), .SE(1'b0), 
      .GCK(n_122_1));
   DFF_X1 \values_reg[98][15]  (.D(values[15]), .CK(n_122_1), .Q(
      \values[98] [15]), .QN());
   DFF_X1 \values_reg[98][14]  (.D(values[14]), .CK(n_122_1), .Q(
      \values[98] [14]), .QN());
   DFF_X1 \values_reg[98][13]  (.D(values[13]), .CK(n_122_1), .Q(
      \values[98] [13]), .QN());
   DFF_X1 \values_reg[98][12]  (.D(values[12]), .CK(n_122_1), .Q(
      \values[98] [12]), .QN());
   DFF_X1 \values_reg[98][11]  (.D(values[11]), .CK(n_122_1), .Q(
      \values[98] [11]), .QN());
   DFF_X1 \values_reg[98][10]  (.D(values[10]), .CK(n_122_1), .Q(
      \values[98] [10]), .QN());
   DFF_X1 \values_reg[98][9]  (.D(values[9]), .CK(n_122_1), .Q(\values[98] [9]), 
      .QN());
   DFF_X1 \values_reg[98][8]  (.D(values[8]), .CK(n_122_1), .Q(\values[98] [8]), 
      .QN());
   DFF_X1 \values_reg[98][7]  (.D(values[7]), .CK(n_122_1), .Q(\values[98] [7]), 
      .QN());
   DFF_X1 \values_reg[98][6]  (.D(values[6]), .CK(n_122_1), .Q(\values[98] [6]), 
      .QN());
   DFF_X1 \values_reg[98][5]  (.D(values[5]), .CK(n_122_1), .Q(\values[98] [5]), 
      .QN());
   DFF_X1 \values_reg[98][4]  (.D(values[4]), .CK(n_122_1), .Q(\values[98] [4]), 
      .QN());
   DFF_X1 \values_reg[98][3]  (.D(values[3]), .CK(n_122_1), .Q(\values[98] [3]), 
      .QN());
   DFF_X1 \values_reg[98][2]  (.D(values[2]), .CK(n_122_1), .Q(\values[98] [2]), 
      .QN());
   DFF_X1 \values_reg[98][1]  (.D(values[1]), .CK(n_122_1), .Q(\values[98] [1]), 
      .QN());
   DFF_X1 \values_reg[98][0]  (.D(values[0]), .CK(n_122_1), .Q(\values[98] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[99]_reg  (.CK(clk), .E(n_99), .SE(1'b0), 
      .GCK(n_122_2));
   DFF_X1 \values_reg[99][15]  (.D(values[15]), .CK(n_122_2), .Q(
      \values[99] [15]), .QN());
   DFF_X1 \values_reg[99][14]  (.D(values[14]), .CK(n_122_2), .Q(
      \values[99] [14]), .QN());
   DFF_X1 \values_reg[99][13]  (.D(values[13]), .CK(n_122_2), .Q(
      \values[99] [13]), .QN());
   DFF_X1 \values_reg[99][12]  (.D(values[12]), .CK(n_122_2), .Q(
      \values[99] [12]), .QN());
   DFF_X1 \values_reg[99][11]  (.D(values[11]), .CK(n_122_2), .Q(
      \values[99] [11]), .QN());
   DFF_X1 \values_reg[99][10]  (.D(values[10]), .CK(n_122_2), .Q(
      \values[99] [10]), .QN());
   DFF_X1 \values_reg[99][9]  (.D(values[9]), .CK(n_122_2), .Q(\values[99] [9]), 
      .QN());
   DFF_X1 \values_reg[99][8]  (.D(values[8]), .CK(n_122_2), .Q(\values[99] [8]), 
      .QN());
   DFF_X1 \values_reg[99][7]  (.D(values[7]), .CK(n_122_2), .Q(\values[99] [7]), 
      .QN());
   DFF_X1 \values_reg[99][6]  (.D(values[6]), .CK(n_122_2), .Q(\values[99] [6]), 
      .QN());
   DFF_X1 \values_reg[99][5]  (.D(values[5]), .CK(n_122_2), .Q(\values[99] [5]), 
      .QN());
   DFF_X1 \values_reg[99][4]  (.D(values[4]), .CK(n_122_2), .Q(\values[99] [4]), 
      .QN());
   DFF_X1 \values_reg[99][3]  (.D(values[3]), .CK(n_122_2), .Q(\values[99] [3]), 
      .QN());
   DFF_X1 \values_reg[99][2]  (.D(values[2]), .CK(n_122_2), .Q(\values[99] [2]), 
      .QN());
   DFF_X1 \values_reg[99][1]  (.D(values[1]), .CK(n_122_2), .Q(\values[99] [1]), 
      .QN());
   DFF_X1 \values_reg[99][0]  (.D(values[0]), .CK(n_122_2), .Q(\values[99] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[100]_reg  (.CK(clk), .E(n_100), .SE(1'b0), 
      .GCK(n_122_3));
   DFF_X1 \values_reg[100][15]  (.D(values[15]), .CK(n_122_3), .Q(
      \values[100] [15]), .QN());
   DFF_X1 \values_reg[100][14]  (.D(values[14]), .CK(n_122_3), .Q(
      \values[100] [14]), .QN());
   DFF_X1 \values_reg[100][13]  (.D(values[13]), .CK(n_122_3), .Q(
      \values[100] [13]), .QN());
   DFF_X1 \values_reg[100][12]  (.D(values[12]), .CK(n_122_3), .Q(
      \values[100] [12]), .QN());
   DFF_X1 \values_reg[100][11]  (.D(values[11]), .CK(n_122_3), .Q(
      \values[100] [11]), .QN());
   DFF_X1 \values_reg[100][10]  (.D(values[10]), .CK(n_122_3), .Q(
      \values[100] [10]), .QN());
   DFF_X1 \values_reg[100][9]  (.D(values[9]), .CK(n_122_3), .Q(\values[100] [9]), 
      .QN());
   DFF_X1 \values_reg[100][8]  (.D(values[8]), .CK(n_122_3), .Q(\values[100] [8]), 
      .QN());
   DFF_X1 \values_reg[100][7]  (.D(values[7]), .CK(n_122_3), .Q(\values[100] [7]), 
      .QN());
   DFF_X1 \values_reg[100][6]  (.D(values[6]), .CK(n_122_3), .Q(\values[100] [6]), 
      .QN());
   DFF_X1 \values_reg[100][5]  (.D(values[5]), .CK(n_122_3), .Q(\values[100] [5]), 
      .QN());
   DFF_X1 \values_reg[100][4]  (.D(values[4]), .CK(n_122_3), .Q(\values[100] [4]), 
      .QN());
   DFF_X1 \values_reg[100][3]  (.D(values[3]), .CK(n_122_3), .Q(\values[100] [3]), 
      .QN());
   DFF_X1 \values_reg[100][2]  (.D(values[2]), .CK(n_122_3), .Q(\values[100] [2]), 
      .QN());
   DFF_X1 \values_reg[100][1]  (.D(values[1]), .CK(n_122_3), .Q(\values[100] [1]), 
      .QN());
   DFF_X1 \values_reg[100][0]  (.D(values[0]), .CK(n_122_3), .Q(\values[100] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[101]_reg  (.CK(clk), .E(n_101), .SE(1'b0), 
      .GCK(n_122_4));
   DFF_X1 \values_reg[101][15]  (.D(values[15]), .CK(n_122_4), .Q(
      \values[101] [15]), .QN());
   DFF_X1 \values_reg[101][14]  (.D(values[14]), .CK(n_122_4), .Q(
      \values[101] [14]), .QN());
   DFF_X1 \values_reg[101][13]  (.D(values[13]), .CK(n_122_4), .Q(
      \values[101] [13]), .QN());
   DFF_X1 \values_reg[101][12]  (.D(values[12]), .CK(n_122_4), .Q(
      \values[101] [12]), .QN());
   DFF_X1 \values_reg[101][11]  (.D(values[11]), .CK(n_122_4), .Q(
      \values[101] [11]), .QN());
   DFF_X1 \values_reg[101][10]  (.D(values[10]), .CK(n_122_4), .Q(
      \values[101] [10]), .QN());
   DFF_X1 \values_reg[101][9]  (.D(values[9]), .CK(n_122_4), .Q(\values[101] [9]), 
      .QN());
   DFF_X1 \values_reg[101][8]  (.D(values[8]), .CK(n_122_4), .Q(\values[101] [8]), 
      .QN());
   DFF_X1 \values_reg[101][7]  (.D(values[7]), .CK(n_122_4), .Q(\values[101] [7]), 
      .QN());
   DFF_X1 \values_reg[101][6]  (.D(values[6]), .CK(n_122_4), .Q(\values[101] [6]), 
      .QN());
   DFF_X1 \values_reg[101][5]  (.D(values[5]), .CK(n_122_4), .Q(\values[101] [5]), 
      .QN());
   DFF_X1 \values_reg[101][4]  (.D(values[4]), .CK(n_122_4), .Q(\values[101] [4]), 
      .QN());
   DFF_X1 \values_reg[101][3]  (.D(values[3]), .CK(n_122_4), .Q(\values[101] [3]), 
      .QN());
   DFF_X1 \values_reg[101][2]  (.D(values[2]), .CK(n_122_4), .Q(\values[101] [2]), 
      .QN());
   DFF_X1 \values_reg[101][1]  (.D(values[1]), .CK(n_122_4), .Q(\values[101] [1]), 
      .QN());
   DFF_X1 \values_reg[101][0]  (.D(values[0]), .CK(n_122_4), .Q(\values[101] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[102]_reg  (.CK(clk), .E(n_102), .SE(1'b0), 
      .GCK(n_122_5));
   DFF_X1 \values_reg[102][15]  (.D(values[15]), .CK(n_122_5), .Q(
      \values[102] [15]), .QN());
   DFF_X1 \values_reg[102][14]  (.D(values[14]), .CK(n_122_5), .Q(
      \values[102] [14]), .QN());
   DFF_X1 \values_reg[102][13]  (.D(values[13]), .CK(n_122_5), .Q(
      \values[102] [13]), .QN());
   DFF_X1 \values_reg[102][12]  (.D(values[12]), .CK(n_122_5), .Q(
      \values[102] [12]), .QN());
   DFF_X1 \values_reg[102][11]  (.D(values[11]), .CK(n_122_5), .Q(
      \values[102] [11]), .QN());
   DFF_X1 \values_reg[102][10]  (.D(values[10]), .CK(n_122_5), .Q(
      \values[102] [10]), .QN());
   DFF_X1 \values_reg[102][9]  (.D(values[9]), .CK(n_122_5), .Q(\values[102] [9]), 
      .QN());
   DFF_X1 \values_reg[102][8]  (.D(values[8]), .CK(n_122_5), .Q(\values[102] [8]), 
      .QN());
   DFF_X1 \values_reg[102][7]  (.D(values[7]), .CK(n_122_5), .Q(\values[102] [7]), 
      .QN());
   DFF_X1 \values_reg[102][6]  (.D(values[6]), .CK(n_122_5), .Q(\values[102] [6]), 
      .QN());
   DFF_X1 \values_reg[102][5]  (.D(values[5]), .CK(n_122_5), .Q(\values[102] [5]), 
      .QN());
   DFF_X1 \values_reg[102][4]  (.D(values[4]), .CK(n_122_5), .Q(\values[102] [4]), 
      .QN());
   DFF_X1 \values_reg[102][3]  (.D(values[3]), .CK(n_122_5), .Q(\values[102] [3]), 
      .QN());
   DFF_X1 \values_reg[102][2]  (.D(values[2]), .CK(n_122_5), .Q(\values[102] [2]), 
      .QN());
   DFF_X1 \values_reg[102][1]  (.D(values[1]), .CK(n_122_5), .Q(\values[102] [1]), 
      .QN());
   DFF_X1 \values_reg[102][0]  (.D(values[0]), .CK(n_122_5), .Q(\values[102] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[103]_reg  (.CK(clk), .E(n_103), .SE(1'b0), 
      .GCK(n_122_6));
   DFF_X1 \values_reg[103][15]  (.D(values[15]), .CK(n_122_6), .Q(
      \values[103] [15]), .QN());
   DFF_X1 \values_reg[103][14]  (.D(values[14]), .CK(n_122_6), .Q(
      \values[103] [14]), .QN());
   DFF_X1 \values_reg[103][13]  (.D(values[13]), .CK(n_122_6), .Q(
      \values[103] [13]), .QN());
   DFF_X1 \values_reg[103][12]  (.D(values[12]), .CK(n_122_6), .Q(
      \values[103] [12]), .QN());
   DFF_X1 \values_reg[103][11]  (.D(values[11]), .CK(n_122_6), .Q(
      \values[103] [11]), .QN());
   DFF_X1 \values_reg[103][10]  (.D(values[10]), .CK(n_122_6), .Q(
      \values[103] [10]), .QN());
   DFF_X1 \values_reg[103][9]  (.D(values[9]), .CK(n_122_6), .Q(\values[103] [9]), 
      .QN());
   DFF_X1 \values_reg[103][8]  (.D(values[8]), .CK(n_122_6), .Q(\values[103] [8]), 
      .QN());
   DFF_X1 \values_reg[103][7]  (.D(values[7]), .CK(n_122_6), .Q(\values[103] [7]), 
      .QN());
   DFF_X1 \values_reg[103][6]  (.D(values[6]), .CK(n_122_6), .Q(\values[103] [6]), 
      .QN());
   DFF_X1 \values_reg[103][5]  (.D(values[5]), .CK(n_122_6), .Q(\values[103] [5]), 
      .QN());
   DFF_X1 \values_reg[103][4]  (.D(values[4]), .CK(n_122_6), .Q(\values[103] [4]), 
      .QN());
   DFF_X1 \values_reg[103][3]  (.D(values[3]), .CK(n_122_6), .Q(\values[103] [3]), 
      .QN());
   DFF_X1 \values_reg[103][2]  (.D(values[2]), .CK(n_122_6), .Q(\values[103] [2]), 
      .QN());
   DFF_X1 \values_reg[103][1]  (.D(values[1]), .CK(n_122_6), .Q(\values[103] [1]), 
      .QN());
   DFF_X1 \values_reg[103][0]  (.D(values[0]), .CK(n_122_6), .Q(\values[103] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[104]_reg  (.CK(clk), .E(n_104), .SE(1'b0), 
      .GCK(n_122_7));
   DFF_X1 \values_reg[104][15]  (.D(values[15]), .CK(n_122_7), .Q(
      \values[104] [15]), .QN());
   DFF_X1 \values_reg[104][14]  (.D(values[14]), .CK(n_122_7), .Q(
      \values[104] [14]), .QN());
   DFF_X1 \values_reg[104][13]  (.D(values[13]), .CK(n_122_7), .Q(
      \values[104] [13]), .QN());
   DFF_X1 \values_reg[104][12]  (.D(values[12]), .CK(n_122_7), .Q(
      \values[104] [12]), .QN());
   DFF_X1 \values_reg[104][11]  (.D(values[11]), .CK(n_122_7), .Q(
      \values[104] [11]), .QN());
   DFF_X1 \values_reg[104][10]  (.D(values[10]), .CK(n_122_7), .Q(
      \values[104] [10]), .QN());
   DFF_X1 \values_reg[104][9]  (.D(values[9]), .CK(n_122_7), .Q(\values[104] [9]), 
      .QN());
   DFF_X1 \values_reg[104][8]  (.D(values[8]), .CK(n_122_7), .Q(\values[104] [8]), 
      .QN());
   DFF_X1 \values_reg[104][7]  (.D(values[7]), .CK(n_122_7), .Q(\values[104] [7]), 
      .QN());
   DFF_X1 \values_reg[104][6]  (.D(values[6]), .CK(n_122_7), .Q(\values[104] [6]), 
      .QN());
   DFF_X1 \values_reg[104][5]  (.D(values[5]), .CK(n_122_7), .Q(\values[104] [5]), 
      .QN());
   DFF_X1 \values_reg[104][4]  (.D(values[4]), .CK(n_122_7), .Q(\values[104] [4]), 
      .QN());
   DFF_X1 \values_reg[104][3]  (.D(values[3]), .CK(n_122_7), .Q(\values[104] [3]), 
      .QN());
   DFF_X1 \values_reg[104][2]  (.D(values[2]), .CK(n_122_7), .Q(\values[104] [2]), 
      .QN());
   DFF_X1 \values_reg[104][1]  (.D(values[1]), .CK(n_122_7), .Q(\values[104] [1]), 
      .QN());
   DFF_X1 \values_reg[104][0]  (.D(values[0]), .CK(n_122_7), .Q(\values[104] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[105]_reg  (.CK(clk), .E(n_105), .SE(1'b0), 
      .GCK(n_122_8));
   DFF_X1 \values_reg[105][15]  (.D(values[15]), .CK(n_122_8), .Q(
      \values[105] [15]), .QN());
   DFF_X1 \values_reg[105][14]  (.D(values[14]), .CK(n_122_8), .Q(
      \values[105] [14]), .QN());
   DFF_X1 \values_reg[105][13]  (.D(values[13]), .CK(n_122_8), .Q(
      \values[105] [13]), .QN());
   DFF_X1 \values_reg[105][12]  (.D(values[12]), .CK(n_122_8), .Q(
      \values[105] [12]), .QN());
   DFF_X1 \values_reg[105][11]  (.D(values[11]), .CK(n_122_8), .Q(
      \values[105] [11]), .QN());
   DFF_X1 \values_reg[105][10]  (.D(values[10]), .CK(n_122_8), .Q(
      \values[105] [10]), .QN());
   DFF_X1 \values_reg[105][9]  (.D(values[9]), .CK(n_122_8), .Q(\values[105] [9]), 
      .QN());
   DFF_X1 \values_reg[105][8]  (.D(values[8]), .CK(n_122_8), .Q(\values[105] [8]), 
      .QN());
   DFF_X1 \values_reg[105][7]  (.D(values[7]), .CK(n_122_8), .Q(\values[105] [7]), 
      .QN());
   DFF_X1 \values_reg[105][6]  (.D(values[6]), .CK(n_122_8), .Q(\values[105] [6]), 
      .QN());
   DFF_X1 \values_reg[105][5]  (.D(values[5]), .CK(n_122_8), .Q(\values[105] [5]), 
      .QN());
   DFF_X1 \values_reg[105][4]  (.D(values[4]), .CK(n_122_8), .Q(\values[105] [4]), 
      .QN());
   DFF_X1 \values_reg[105][3]  (.D(values[3]), .CK(n_122_8), .Q(\values[105] [3]), 
      .QN());
   DFF_X1 \values_reg[105][2]  (.D(values[2]), .CK(n_122_8), .Q(\values[105] [2]), 
      .QN());
   DFF_X1 \values_reg[105][1]  (.D(values[1]), .CK(n_122_8), .Q(\values[105] [1]), 
      .QN());
   DFF_X1 \values_reg[105][0]  (.D(values[0]), .CK(n_122_8), .Q(\values[105] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[106]_reg  (.CK(clk), .E(n_106), .SE(1'b0), 
      .GCK(n_122_9));
   DFF_X1 \values_reg[106][15]  (.D(values[15]), .CK(n_122_9), .Q(
      \values[106] [15]), .QN());
   DFF_X1 \values_reg[106][14]  (.D(values[14]), .CK(n_122_9), .Q(
      \values[106] [14]), .QN());
   DFF_X1 \values_reg[106][13]  (.D(values[13]), .CK(n_122_9), .Q(
      \values[106] [13]), .QN());
   DFF_X1 \values_reg[106][12]  (.D(values[12]), .CK(n_122_9), .Q(
      \values[106] [12]), .QN());
   DFF_X1 \values_reg[106][11]  (.D(values[11]), .CK(n_122_9), .Q(
      \values[106] [11]), .QN());
   DFF_X1 \values_reg[106][10]  (.D(values[10]), .CK(n_122_9), .Q(
      \values[106] [10]), .QN());
   DFF_X1 \values_reg[106][9]  (.D(values[9]), .CK(n_122_9), .Q(\values[106] [9]), 
      .QN());
   DFF_X1 \values_reg[106][8]  (.D(values[8]), .CK(n_122_9), .Q(\values[106] [8]), 
      .QN());
   DFF_X1 \values_reg[106][7]  (.D(values[7]), .CK(n_122_9), .Q(\values[106] [7]), 
      .QN());
   DFF_X1 \values_reg[106][6]  (.D(values[6]), .CK(n_122_9), .Q(\values[106] [6]), 
      .QN());
   DFF_X1 \values_reg[106][5]  (.D(values[5]), .CK(n_122_9), .Q(\values[106] [5]), 
      .QN());
   DFF_X1 \values_reg[106][4]  (.D(values[4]), .CK(n_122_9), .Q(\values[106] [4]), 
      .QN());
   DFF_X1 \values_reg[106][3]  (.D(values[3]), .CK(n_122_9), .Q(\values[106] [3]), 
      .QN());
   DFF_X1 \values_reg[106][2]  (.D(values[2]), .CK(n_122_9), .Q(\values[106] [2]), 
      .QN());
   DFF_X1 \values_reg[106][1]  (.D(values[1]), .CK(n_122_9), .Q(\values[106] [1]), 
      .QN());
   DFF_X1 \values_reg[106][0]  (.D(values[0]), .CK(n_122_9), .Q(\values[106] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[107]_reg  (.CK(clk), .E(n_107), .SE(1'b0), 
      .GCK(n_122_10));
   DFF_X1 \values_reg[107][15]  (.D(values[15]), .CK(n_122_10), .Q(
      \values[107] [15]), .QN());
   DFF_X1 \values_reg[107][14]  (.D(values[14]), .CK(n_122_10), .Q(
      \values[107] [14]), .QN());
   DFF_X1 \values_reg[107][13]  (.D(values[13]), .CK(n_122_10), .Q(
      \values[107] [13]), .QN());
   DFF_X1 \values_reg[107][12]  (.D(values[12]), .CK(n_122_10), .Q(
      \values[107] [12]), .QN());
   DFF_X1 \values_reg[107][11]  (.D(values[11]), .CK(n_122_10), .Q(
      \values[107] [11]), .QN());
   DFF_X1 \values_reg[107][10]  (.D(values[10]), .CK(n_122_10), .Q(
      \values[107] [10]), .QN());
   DFF_X1 \values_reg[107][9]  (.D(values[9]), .CK(n_122_10), .Q(
      \values[107] [9]), .QN());
   DFF_X1 \values_reg[107][8]  (.D(values[8]), .CK(n_122_10), .Q(
      \values[107] [8]), .QN());
   DFF_X1 \values_reg[107][7]  (.D(values[7]), .CK(n_122_10), .Q(
      \values[107] [7]), .QN());
   DFF_X1 \values_reg[107][6]  (.D(values[6]), .CK(n_122_10), .Q(
      \values[107] [6]), .QN());
   DFF_X1 \values_reg[107][5]  (.D(values[5]), .CK(n_122_10), .Q(
      \values[107] [5]), .QN());
   DFF_X1 \values_reg[107][4]  (.D(values[4]), .CK(n_122_10), .Q(
      \values[107] [4]), .QN());
   DFF_X1 \values_reg[107][3]  (.D(values[3]), .CK(n_122_10), .Q(
      \values[107] [3]), .QN());
   DFF_X1 \values_reg[107][2]  (.D(values[2]), .CK(n_122_10), .Q(
      \values[107] [2]), .QN());
   DFF_X1 \values_reg[107][1]  (.D(values[1]), .CK(n_122_10), .Q(
      \values[107] [1]), .QN());
   DFF_X1 \values_reg[107][0]  (.D(values[0]), .CK(n_122_10), .Q(
      \values[107] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[108]_reg  (.CK(clk), .E(n_108), .SE(1'b0), 
      .GCK(n_122_11));
   DFF_X1 \values_reg[108][15]  (.D(values[15]), .CK(n_122_11), .Q(
      \values[108] [15]), .QN());
   DFF_X1 \values_reg[108][14]  (.D(values[14]), .CK(n_122_11), .Q(
      \values[108] [14]), .QN());
   DFF_X1 \values_reg[108][13]  (.D(values[13]), .CK(n_122_11), .Q(
      \values[108] [13]), .QN());
   DFF_X1 \values_reg[108][12]  (.D(values[12]), .CK(n_122_11), .Q(
      \values[108] [12]), .QN());
   DFF_X1 \values_reg[108][11]  (.D(values[11]), .CK(n_122_11), .Q(
      \values[108] [11]), .QN());
   DFF_X1 \values_reg[108][10]  (.D(values[10]), .CK(n_122_11), .Q(
      \values[108] [10]), .QN());
   DFF_X1 \values_reg[108][9]  (.D(values[9]), .CK(n_122_11), .Q(
      \values[108] [9]), .QN());
   DFF_X1 \values_reg[108][8]  (.D(values[8]), .CK(n_122_11), .Q(
      \values[108] [8]), .QN());
   DFF_X1 \values_reg[108][7]  (.D(values[7]), .CK(n_122_11), .Q(
      \values[108] [7]), .QN());
   DFF_X1 \values_reg[108][6]  (.D(values[6]), .CK(n_122_11), .Q(
      \values[108] [6]), .QN());
   DFF_X1 \values_reg[108][5]  (.D(values[5]), .CK(n_122_11), .Q(
      \values[108] [5]), .QN());
   DFF_X1 \values_reg[108][4]  (.D(values[4]), .CK(n_122_11), .Q(
      \values[108] [4]), .QN());
   DFF_X1 \values_reg[108][3]  (.D(values[3]), .CK(n_122_11), .Q(
      \values[108] [3]), .QN());
   DFF_X1 \values_reg[108][2]  (.D(values[2]), .CK(n_122_11), .Q(
      \values[108] [2]), .QN());
   DFF_X1 \values_reg[108][1]  (.D(values[1]), .CK(n_122_11), .Q(
      \values[108] [1]), .QN());
   DFF_X1 \values_reg[108][0]  (.D(values[0]), .CK(n_122_11), .Q(
      \values[108] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[109]_reg  (.CK(clk), .E(n_109), .SE(1'b0), 
      .GCK(n_122_12));
   DFF_X1 \values_reg[109][15]  (.D(values[15]), .CK(n_122_12), .Q(
      \values[109] [15]), .QN());
   DFF_X1 \values_reg[109][14]  (.D(values[14]), .CK(n_122_12), .Q(
      \values[109] [14]), .QN());
   DFF_X1 \values_reg[109][13]  (.D(values[13]), .CK(n_122_12), .Q(
      \values[109] [13]), .QN());
   DFF_X1 \values_reg[109][12]  (.D(values[12]), .CK(n_122_12), .Q(
      \values[109] [12]), .QN());
   DFF_X1 \values_reg[109][11]  (.D(values[11]), .CK(n_122_12), .Q(
      \values[109] [11]), .QN());
   DFF_X1 \values_reg[109][10]  (.D(values[10]), .CK(n_122_12), .Q(
      \values[109] [10]), .QN());
   DFF_X1 \values_reg[109][9]  (.D(values[9]), .CK(n_122_12), .Q(
      \values[109] [9]), .QN());
   DFF_X1 \values_reg[109][8]  (.D(values[8]), .CK(n_122_12), .Q(
      \values[109] [8]), .QN());
   DFF_X1 \values_reg[109][7]  (.D(values[7]), .CK(n_122_12), .Q(
      \values[109] [7]), .QN());
   DFF_X1 \values_reg[109][6]  (.D(values[6]), .CK(n_122_12), .Q(
      \values[109] [6]), .QN());
   DFF_X1 \values_reg[109][5]  (.D(values[5]), .CK(n_122_12), .Q(
      \values[109] [5]), .QN());
   DFF_X1 \values_reg[109][4]  (.D(values[4]), .CK(n_122_12), .Q(
      \values[109] [4]), .QN());
   DFF_X1 \values_reg[109][3]  (.D(values[3]), .CK(n_122_12), .Q(
      \values[109] [3]), .QN());
   DFF_X1 \values_reg[109][2]  (.D(values[2]), .CK(n_122_12), .Q(
      \values[109] [2]), .QN());
   DFF_X1 \values_reg[109][1]  (.D(values[1]), .CK(n_122_12), .Q(
      \values[109] [1]), .QN());
   DFF_X1 \values_reg[109][0]  (.D(values[0]), .CK(n_122_12), .Q(
      \values[109] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[110]_reg  (.CK(clk), .E(n_110), .SE(1'b0), 
      .GCK(n_122_13));
   DFF_X1 \values_reg[110][15]  (.D(values[15]), .CK(n_122_13), .Q(
      \values[110] [15]), .QN());
   DFF_X1 \values_reg[110][14]  (.D(values[14]), .CK(n_122_13), .Q(
      \values[110] [14]), .QN());
   DFF_X1 \values_reg[110][13]  (.D(values[13]), .CK(n_122_13), .Q(
      \values[110] [13]), .QN());
   DFF_X1 \values_reg[110][12]  (.D(values[12]), .CK(n_122_13), .Q(
      \values[110] [12]), .QN());
   DFF_X1 \values_reg[110][11]  (.D(values[11]), .CK(n_122_13), .Q(
      \values[110] [11]), .QN());
   DFF_X1 \values_reg[110][10]  (.D(values[10]), .CK(n_122_13), .Q(
      \values[110] [10]), .QN());
   DFF_X1 \values_reg[110][9]  (.D(values[9]), .CK(n_122_13), .Q(
      \values[110] [9]), .QN());
   DFF_X1 \values_reg[110][8]  (.D(values[8]), .CK(n_122_13), .Q(
      \values[110] [8]), .QN());
   DFF_X1 \values_reg[110][7]  (.D(values[7]), .CK(n_122_13), .Q(
      \values[110] [7]), .QN());
   DFF_X1 \values_reg[110][6]  (.D(values[6]), .CK(n_122_13), .Q(
      \values[110] [6]), .QN());
   DFF_X1 \values_reg[110][5]  (.D(values[5]), .CK(n_122_13), .Q(
      \values[110] [5]), .QN());
   DFF_X1 \values_reg[110][4]  (.D(values[4]), .CK(n_122_13), .Q(
      \values[110] [4]), .QN());
   DFF_X1 \values_reg[110][3]  (.D(values[3]), .CK(n_122_13), .Q(
      \values[110] [3]), .QN());
   DFF_X1 \values_reg[110][2]  (.D(values[2]), .CK(n_122_13), .Q(
      \values[110] [2]), .QN());
   DFF_X1 \values_reg[110][1]  (.D(values[1]), .CK(n_122_13), .Q(
      \values[110] [1]), .QN());
   DFF_X1 \values_reg[110][0]  (.D(values[0]), .CK(n_122_13), .Q(
      \values[110] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[111]_reg  (.CK(clk), .E(n_111), .SE(1'b0), 
      .GCK(n_122_14));
   DFF_X1 \values_reg[111][15]  (.D(values[15]), .CK(n_122_14), .Q(
      \values[111] [15]), .QN());
   DFF_X1 \values_reg[111][14]  (.D(values[14]), .CK(n_122_14), .Q(
      \values[111] [14]), .QN());
   DFF_X1 \values_reg[111][13]  (.D(values[13]), .CK(n_122_14), .Q(
      \values[111] [13]), .QN());
   DFF_X1 \values_reg[111][12]  (.D(values[12]), .CK(n_122_14), .Q(
      \values[111] [12]), .QN());
   DFF_X1 \values_reg[111][11]  (.D(values[11]), .CK(n_122_14), .Q(
      \values[111] [11]), .QN());
   DFF_X1 \values_reg[111][10]  (.D(values[10]), .CK(n_122_14), .Q(
      \values[111] [10]), .QN());
   DFF_X1 \values_reg[111][9]  (.D(values[9]), .CK(n_122_14), .Q(
      \values[111] [9]), .QN());
   DFF_X1 \values_reg[111][8]  (.D(values[8]), .CK(n_122_14), .Q(
      \values[111] [8]), .QN());
   DFF_X1 \values_reg[111][7]  (.D(values[7]), .CK(n_122_14), .Q(
      \values[111] [7]), .QN());
   DFF_X1 \values_reg[111][6]  (.D(values[6]), .CK(n_122_14), .Q(
      \values[111] [6]), .QN());
   DFF_X1 \values_reg[111][5]  (.D(values[5]), .CK(n_122_14), .Q(
      \values[111] [5]), .QN());
   DFF_X1 \values_reg[111][4]  (.D(values[4]), .CK(n_122_14), .Q(
      \values[111] [4]), .QN());
   DFF_X1 \values_reg[111][3]  (.D(values[3]), .CK(n_122_14), .Q(
      \values[111] [3]), .QN());
   DFF_X1 \values_reg[111][2]  (.D(values[2]), .CK(n_122_14), .Q(
      \values[111] [2]), .QN());
   DFF_X1 \values_reg[111][1]  (.D(values[1]), .CK(n_122_14), .Q(
      \values[111] [1]), .QN());
   DFF_X1 \values_reg[111][0]  (.D(values[0]), .CK(n_122_14), .Q(
      \values[111] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[112]_reg  (.CK(clk), .E(n_112), .SE(1'b0), 
      .GCK(n_122_15));
   DFF_X1 \values_reg[112][15]  (.D(values[15]), .CK(n_122_15), .Q(
      \values[112] [15]), .QN());
   DFF_X1 \values_reg[112][14]  (.D(values[14]), .CK(n_122_15), .Q(
      \values[112] [14]), .QN());
   DFF_X1 \values_reg[112][13]  (.D(values[13]), .CK(n_122_15), .Q(
      \values[112] [13]), .QN());
   DFF_X1 \values_reg[112][12]  (.D(values[12]), .CK(n_122_15), .Q(
      \values[112] [12]), .QN());
   DFF_X1 \values_reg[112][11]  (.D(values[11]), .CK(n_122_15), .Q(
      \values[112] [11]), .QN());
   DFF_X1 \values_reg[112][10]  (.D(values[10]), .CK(n_122_15), .Q(
      \values[112] [10]), .QN());
   DFF_X1 \values_reg[112][9]  (.D(values[9]), .CK(n_122_15), .Q(
      \values[112] [9]), .QN());
   DFF_X1 \values_reg[112][8]  (.D(values[8]), .CK(n_122_15), .Q(
      \values[112] [8]), .QN());
   DFF_X1 \values_reg[112][7]  (.D(values[7]), .CK(n_122_15), .Q(
      \values[112] [7]), .QN());
   DFF_X1 \values_reg[112][6]  (.D(values[6]), .CK(n_122_15), .Q(
      \values[112] [6]), .QN());
   DFF_X1 \values_reg[112][5]  (.D(values[5]), .CK(n_122_15), .Q(
      \values[112] [5]), .QN());
   DFF_X1 \values_reg[112][4]  (.D(values[4]), .CK(n_122_15), .Q(
      \values[112] [4]), .QN());
   DFF_X1 \values_reg[112][3]  (.D(values[3]), .CK(n_122_15), .Q(
      \values[112] [3]), .QN());
   DFF_X1 \values_reg[112][2]  (.D(values[2]), .CK(n_122_15), .Q(
      \values[112] [2]), .QN());
   DFF_X1 \values_reg[112][1]  (.D(values[1]), .CK(n_122_15), .Q(
      \values[112] [1]), .QN());
   DFF_X1 \values_reg[112][0]  (.D(values[0]), .CK(n_122_15), .Q(
      \values[112] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[113]_reg  (.CK(clk), .E(n_113), .SE(1'b0), 
      .GCK(n_122_16));
   DFF_X1 \values_reg[113][15]  (.D(values[15]), .CK(n_122_16), .Q(
      \values[113] [15]), .QN());
   DFF_X1 \values_reg[113][14]  (.D(values[14]), .CK(n_122_16), .Q(
      \values[113] [14]), .QN());
   DFF_X1 \values_reg[113][13]  (.D(values[13]), .CK(n_122_16), .Q(
      \values[113] [13]), .QN());
   DFF_X1 \values_reg[113][12]  (.D(values[12]), .CK(n_122_16), .Q(
      \values[113] [12]), .QN());
   DFF_X1 \values_reg[113][11]  (.D(values[11]), .CK(n_122_16), .Q(
      \values[113] [11]), .QN());
   DFF_X1 \values_reg[113][10]  (.D(values[10]), .CK(n_122_16), .Q(
      \values[113] [10]), .QN());
   DFF_X1 \values_reg[113][9]  (.D(values[9]), .CK(n_122_16), .Q(
      \values[113] [9]), .QN());
   DFF_X1 \values_reg[113][8]  (.D(values[8]), .CK(n_122_16), .Q(
      \values[113] [8]), .QN());
   DFF_X1 \values_reg[113][7]  (.D(values[7]), .CK(n_122_16), .Q(
      \values[113] [7]), .QN());
   DFF_X1 \values_reg[113][6]  (.D(values[6]), .CK(n_122_16), .Q(
      \values[113] [6]), .QN());
   DFF_X1 \values_reg[113][5]  (.D(values[5]), .CK(n_122_16), .Q(
      \values[113] [5]), .QN());
   DFF_X1 \values_reg[113][4]  (.D(values[4]), .CK(n_122_16), .Q(
      \values[113] [4]), .QN());
   DFF_X1 \values_reg[113][3]  (.D(values[3]), .CK(n_122_16), .Q(
      \values[113] [3]), .QN());
   DFF_X1 \values_reg[113][2]  (.D(values[2]), .CK(n_122_16), .Q(
      \values[113] [2]), .QN());
   DFF_X1 \values_reg[113][1]  (.D(values[1]), .CK(n_122_16), .Q(
      \values[113] [1]), .QN());
   DFF_X1 \values_reg[113][0]  (.D(values[0]), .CK(n_122_16), .Q(
      \values[113] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[114]_reg  (.CK(clk), .E(n_114), .SE(1'b0), 
      .GCK(n_122_17));
   DFF_X1 \values_reg[114][15]  (.D(values[15]), .CK(n_122_17), .Q(
      \values[114] [15]), .QN());
   DFF_X1 \values_reg[114][14]  (.D(values[14]), .CK(n_122_17), .Q(
      \values[114] [14]), .QN());
   DFF_X1 \values_reg[114][13]  (.D(values[13]), .CK(n_122_17), .Q(
      \values[114] [13]), .QN());
   DFF_X1 \values_reg[114][12]  (.D(values[12]), .CK(n_122_17), .Q(
      \values[114] [12]), .QN());
   DFF_X1 \values_reg[114][11]  (.D(values[11]), .CK(n_122_17), .Q(
      \values[114] [11]), .QN());
   DFF_X1 \values_reg[114][10]  (.D(values[10]), .CK(n_122_17), .Q(
      \values[114] [10]), .QN());
   DFF_X1 \values_reg[114][9]  (.D(values[9]), .CK(n_122_17), .Q(
      \values[114] [9]), .QN());
   DFF_X1 \values_reg[114][8]  (.D(values[8]), .CK(n_122_17), .Q(
      \values[114] [8]), .QN());
   DFF_X1 \values_reg[114][7]  (.D(values[7]), .CK(n_122_17), .Q(
      \values[114] [7]), .QN());
   DFF_X1 \values_reg[114][6]  (.D(values[6]), .CK(n_122_17), .Q(
      \values[114] [6]), .QN());
   DFF_X1 \values_reg[114][5]  (.D(values[5]), .CK(n_122_17), .Q(
      \values[114] [5]), .QN());
   DFF_X1 \values_reg[114][4]  (.D(values[4]), .CK(n_122_17), .Q(
      \values[114] [4]), .QN());
   DFF_X1 \values_reg[114][3]  (.D(values[3]), .CK(n_122_17), .Q(
      \values[114] [3]), .QN());
   DFF_X1 \values_reg[114][2]  (.D(values[2]), .CK(n_122_17), .Q(
      \values[114] [2]), .QN());
   DFF_X1 \values_reg[114][1]  (.D(values[1]), .CK(n_122_17), .Q(
      \values[114] [1]), .QN());
   DFF_X1 \values_reg[114][0]  (.D(values[0]), .CK(n_122_17), .Q(
      \values[114] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[115]_reg  (.CK(clk), .E(n_115), .SE(1'b0), 
      .GCK(n_122_18));
   DFF_X1 \values_reg[115][15]  (.D(values[15]), .CK(n_122_18), .Q(
      \values[115] [15]), .QN());
   DFF_X1 \values_reg[115][14]  (.D(values[14]), .CK(n_122_18), .Q(
      \values[115] [14]), .QN());
   DFF_X1 \values_reg[115][13]  (.D(values[13]), .CK(n_122_18), .Q(
      \values[115] [13]), .QN());
   DFF_X1 \values_reg[115][12]  (.D(values[12]), .CK(n_122_18), .Q(
      \values[115] [12]), .QN());
   DFF_X1 \values_reg[115][11]  (.D(values[11]), .CK(n_122_18), .Q(
      \values[115] [11]), .QN());
   DFF_X1 \values_reg[115][10]  (.D(values[10]), .CK(n_122_18), .Q(
      \values[115] [10]), .QN());
   DFF_X1 \values_reg[115][9]  (.D(values[9]), .CK(n_122_18), .Q(
      \values[115] [9]), .QN());
   DFF_X1 \values_reg[115][8]  (.D(values[8]), .CK(n_122_18), .Q(
      \values[115] [8]), .QN());
   DFF_X1 \values_reg[115][7]  (.D(values[7]), .CK(n_122_18), .Q(
      \values[115] [7]), .QN());
   DFF_X1 \values_reg[115][6]  (.D(values[6]), .CK(n_122_18), .Q(
      \values[115] [6]), .QN());
   DFF_X1 \values_reg[115][5]  (.D(values[5]), .CK(n_122_18), .Q(
      \values[115] [5]), .QN());
   DFF_X1 \values_reg[115][4]  (.D(values[4]), .CK(n_122_18), .Q(
      \values[115] [4]), .QN());
   DFF_X1 \values_reg[115][3]  (.D(values[3]), .CK(n_122_18), .Q(
      \values[115] [3]), .QN());
   DFF_X1 \values_reg[115][2]  (.D(values[2]), .CK(n_122_18), .Q(
      \values[115] [2]), .QN());
   DFF_X1 \values_reg[115][1]  (.D(values[1]), .CK(n_122_18), .Q(
      \values[115] [1]), .QN());
   DFF_X1 \values_reg[115][0]  (.D(values[0]), .CK(n_122_18), .Q(
      \values[115] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[116]_reg  (.CK(clk), .E(n_116), .SE(1'b0), 
      .GCK(n_122_19));
   DFF_X1 \values_reg[116][15]  (.D(values[15]), .CK(n_122_19), .Q(
      \values[116] [15]), .QN());
   DFF_X1 \values_reg[116][14]  (.D(values[14]), .CK(n_122_19), .Q(
      \values[116] [14]), .QN());
   DFF_X1 \values_reg[116][13]  (.D(values[13]), .CK(n_122_19), .Q(
      \values[116] [13]), .QN());
   DFF_X1 \values_reg[116][12]  (.D(values[12]), .CK(n_122_19), .Q(
      \values[116] [12]), .QN());
   DFF_X1 \values_reg[116][11]  (.D(values[11]), .CK(n_122_19), .Q(
      \values[116] [11]), .QN());
   DFF_X1 \values_reg[116][10]  (.D(values[10]), .CK(n_122_19), .Q(
      \values[116] [10]), .QN());
   DFF_X1 \values_reg[116][9]  (.D(values[9]), .CK(n_122_19), .Q(
      \values[116] [9]), .QN());
   DFF_X1 \values_reg[116][8]  (.D(values[8]), .CK(n_122_19), .Q(
      \values[116] [8]), .QN());
   DFF_X1 \values_reg[116][7]  (.D(values[7]), .CK(n_122_19), .Q(
      \values[116] [7]), .QN());
   DFF_X1 \values_reg[116][6]  (.D(values[6]), .CK(n_122_19), .Q(
      \values[116] [6]), .QN());
   DFF_X1 \values_reg[116][5]  (.D(values[5]), .CK(n_122_19), .Q(
      \values[116] [5]), .QN());
   DFF_X1 \values_reg[116][4]  (.D(values[4]), .CK(n_122_19), .Q(
      \values[116] [4]), .QN());
   DFF_X1 \values_reg[116][3]  (.D(values[3]), .CK(n_122_19), .Q(
      \values[116] [3]), .QN());
   DFF_X1 \values_reg[116][2]  (.D(values[2]), .CK(n_122_19), .Q(
      \values[116] [2]), .QN());
   DFF_X1 \values_reg[116][1]  (.D(values[1]), .CK(n_122_19), .Q(
      \values[116] [1]), .QN());
   DFF_X1 \values_reg[116][0]  (.D(values[0]), .CK(n_122_19), .Q(
      \values[116] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[117]_reg  (.CK(clk), .E(n_117), .SE(1'b0), 
      .GCK(n_122_20));
   DFF_X1 \values_reg[117][15]  (.D(values[15]), .CK(n_122_20), .Q(
      \values[117] [15]), .QN());
   DFF_X1 \values_reg[117][14]  (.D(values[14]), .CK(n_122_20), .Q(
      \values[117] [14]), .QN());
   DFF_X1 \values_reg[117][13]  (.D(values[13]), .CK(n_122_20), .Q(
      \values[117] [13]), .QN());
   DFF_X1 \values_reg[117][12]  (.D(values[12]), .CK(n_122_20), .Q(
      \values[117] [12]), .QN());
   DFF_X1 \values_reg[117][11]  (.D(values[11]), .CK(n_122_20), .Q(
      \values[117] [11]), .QN());
   DFF_X1 \values_reg[117][10]  (.D(values[10]), .CK(n_122_20), .Q(
      \values[117] [10]), .QN());
   DFF_X1 \values_reg[117][9]  (.D(values[9]), .CK(n_122_20), .Q(
      \values[117] [9]), .QN());
   DFF_X1 \values_reg[117][8]  (.D(values[8]), .CK(n_122_20), .Q(
      \values[117] [8]), .QN());
   DFF_X1 \values_reg[117][7]  (.D(values[7]), .CK(n_122_20), .Q(
      \values[117] [7]), .QN());
   DFF_X1 \values_reg[117][6]  (.D(values[6]), .CK(n_122_20), .Q(
      \values[117] [6]), .QN());
   DFF_X1 \values_reg[117][5]  (.D(values[5]), .CK(n_122_20), .Q(
      \values[117] [5]), .QN());
   DFF_X1 \values_reg[117][4]  (.D(values[4]), .CK(n_122_20), .Q(
      \values[117] [4]), .QN());
   DFF_X1 \values_reg[117][3]  (.D(values[3]), .CK(n_122_20), .Q(
      \values[117] [3]), .QN());
   DFF_X1 \values_reg[117][2]  (.D(values[2]), .CK(n_122_20), .Q(
      \values[117] [2]), .QN());
   DFF_X1 \values_reg[117][1]  (.D(values[1]), .CK(n_122_20), .Q(
      \values[117] [1]), .QN());
   DFF_X1 \values_reg[117][0]  (.D(values[0]), .CK(n_122_20), .Q(
      \values[117] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[118]_reg  (.CK(clk), .E(n_118), .SE(1'b0), 
      .GCK(n_122_21));
   DFF_X1 \values_reg[118][15]  (.D(values[15]), .CK(n_122_21), .Q(
      \values[118] [15]), .QN());
   DFF_X1 \values_reg[118][14]  (.D(values[14]), .CK(n_122_21), .Q(
      \values[118] [14]), .QN());
   DFF_X1 \values_reg[118][13]  (.D(values[13]), .CK(n_122_21), .Q(
      \values[118] [13]), .QN());
   DFF_X1 \values_reg[118][12]  (.D(values[12]), .CK(n_122_21), .Q(
      \values[118] [12]), .QN());
   DFF_X1 \values_reg[118][11]  (.D(values[11]), .CK(n_122_21), .Q(
      \values[118] [11]), .QN());
   DFF_X1 \values_reg[118][10]  (.D(values[10]), .CK(n_122_21), .Q(
      \values[118] [10]), .QN());
   DFF_X1 \values_reg[118][9]  (.D(values[9]), .CK(n_122_21), .Q(
      \values[118] [9]), .QN());
   DFF_X1 \values_reg[118][8]  (.D(values[8]), .CK(n_122_21), .Q(
      \values[118] [8]), .QN());
   DFF_X1 \values_reg[118][7]  (.D(values[7]), .CK(n_122_21), .Q(
      \values[118] [7]), .QN());
   DFF_X1 \values_reg[118][6]  (.D(values[6]), .CK(n_122_21), .Q(
      \values[118] [6]), .QN());
   DFF_X1 \values_reg[118][5]  (.D(values[5]), .CK(n_122_21), .Q(
      \values[118] [5]), .QN());
   DFF_X1 \values_reg[118][4]  (.D(values[4]), .CK(n_122_21), .Q(
      \values[118] [4]), .QN());
   DFF_X1 \values_reg[118][3]  (.D(values[3]), .CK(n_122_21), .Q(
      \values[118] [3]), .QN());
   DFF_X1 \values_reg[118][2]  (.D(values[2]), .CK(n_122_21), .Q(
      \values[118] [2]), .QN());
   DFF_X1 \values_reg[118][1]  (.D(values[1]), .CK(n_122_21), .Q(
      \values[118] [1]), .QN());
   DFF_X1 \values_reg[118][0]  (.D(values[0]), .CK(n_122_21), .Q(
      \values[118] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[119]_reg  (.CK(clk), .E(n_119), .SE(1'b0), 
      .GCK(n_122_22));
   DFF_X1 \values_reg[119][15]  (.D(values[15]), .CK(n_122_22), .Q(
      \values[119] [15]), .QN());
   DFF_X1 \values_reg[119][14]  (.D(values[14]), .CK(n_122_22), .Q(
      \values[119] [14]), .QN());
   DFF_X1 \values_reg[119][13]  (.D(values[13]), .CK(n_122_22), .Q(
      \values[119] [13]), .QN());
   DFF_X1 \values_reg[119][12]  (.D(values[12]), .CK(n_122_22), .Q(
      \values[119] [12]), .QN());
   DFF_X1 \values_reg[119][11]  (.D(values[11]), .CK(n_122_22), .Q(
      \values[119] [11]), .QN());
   DFF_X1 \values_reg[119][10]  (.D(values[10]), .CK(n_122_22), .Q(
      \values[119] [10]), .QN());
   DFF_X1 \values_reg[119][9]  (.D(values[9]), .CK(n_122_22), .Q(
      \values[119] [9]), .QN());
   DFF_X1 \values_reg[119][8]  (.D(values[8]), .CK(n_122_22), .Q(
      \values[119] [8]), .QN());
   DFF_X1 \values_reg[119][7]  (.D(values[7]), .CK(n_122_22), .Q(
      \values[119] [7]), .QN());
   DFF_X1 \values_reg[119][6]  (.D(values[6]), .CK(n_122_22), .Q(
      \values[119] [6]), .QN());
   DFF_X1 \values_reg[119][5]  (.D(values[5]), .CK(n_122_22), .Q(
      \values[119] [5]), .QN());
   DFF_X1 \values_reg[119][4]  (.D(values[4]), .CK(n_122_22), .Q(
      \values[119] [4]), .QN());
   DFF_X1 \values_reg[119][3]  (.D(values[3]), .CK(n_122_22), .Q(
      \values[119] [3]), .QN());
   DFF_X1 \values_reg[119][2]  (.D(values[2]), .CK(n_122_22), .Q(
      \values[119] [2]), .QN());
   DFF_X1 \values_reg[119][1]  (.D(values[1]), .CK(n_122_22), .Q(
      \values[119] [1]), .QN());
   DFF_X1 \values_reg[119][0]  (.D(values[0]), .CK(n_122_22), .Q(
      \values[119] [0]), .QN());
   CLKGATETST_X1 \clk_gate_values_reg[2]_reg  (.CK(clk), .E(n_2), .SE(1'b0), 
      .GCK(n_122_23));
   DFF_X1 \values_reg[2][15]  (.D(values[15]), .CK(n_122_23), .Q(\values[2] [15]), 
      .QN());
   DFF_X1 \values_reg[2][14]  (.D(values[14]), .CK(n_122_23), .Q(\values[2] [14]), 
      .QN());
   DFF_X1 \values_reg[2][13]  (.D(values[13]), .CK(n_122_23), .Q(\values[2] [13]), 
      .QN());
   DFF_X1 \values_reg[2][12]  (.D(values[12]), .CK(n_122_23), .Q(\values[2] [12]), 
      .QN());
   DFF_X1 \values_reg[2][11]  (.D(values[11]), .CK(n_122_23), .Q(\values[2] [11]), 
      .QN());
   DFF_X1 \values_reg[2][10]  (.D(values[10]), .CK(n_122_23), .Q(\values[2] [10]), 
      .QN());
   DFF_X1 \values_reg[2][9]  (.D(values[9]), .CK(n_122_23), .Q(\values[2] [9]), 
      .QN());
   DFF_X1 \values_reg[2][8]  (.D(values[8]), .CK(n_122_23), .Q(\values[2] [8]), 
      .QN());
   DFF_X1 \values_reg[2][7]  (.D(values[7]), .CK(n_122_23), .Q(\values[2] [7]), 
      .QN());
   DFF_X1 \values_reg[2][6]  (.D(values[6]), .CK(n_122_23), .Q(\values[2] [6]), 
      .QN());
   DFF_X1 \values_reg[2][5]  (.D(values[5]), .CK(n_122_23), .Q(\values[2] [5]), 
      .QN());
   DFF_X1 \values_reg[2][4]  (.D(values[4]), .CK(n_122_23), .Q(\values[2] [4]), 
      .QN());
   DFF_X1 \values_reg[2][3]  (.D(values[3]), .CK(n_122_23), .Q(\values[2] [3]), 
      .QN());
   DFF_X1 \values_reg[2][2]  (.D(values[2]), .CK(n_122_23), .Q(\values[2] [2]), 
      .QN());
   DFF_X1 \values_reg[2][1]  (.D(values[1]), .CK(n_122_23), .Q(\values[2] [1]), 
      .QN());
   DFF_X1 \values_reg[2][0]  (.D(values[0]), .CK(n_122_23), .Q(\values[2] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[1]_reg  (.CK(clk), .E(n_1), .SE(1'b0), 
      .GCK(n_122_24));
   DFF_X1 \values_reg[1][15]  (.D(values[15]), .CK(n_122_24), .Q(\values[1] [15]), 
      .QN());
   DFF_X1 \values_reg[1][14]  (.D(values[14]), .CK(n_122_24), .Q(\values[1] [14]), 
      .QN());
   DFF_X1 \values_reg[1][13]  (.D(values[13]), .CK(n_122_24), .Q(\values[1] [13]), 
      .QN());
   DFF_X1 \values_reg[1][12]  (.D(values[12]), .CK(n_122_24), .Q(\values[1] [12]), 
      .QN());
   DFF_X1 \values_reg[1][11]  (.D(values[11]), .CK(n_122_24), .Q(\values[1] [11]), 
      .QN());
   DFF_X1 \values_reg[1][10]  (.D(values[10]), .CK(n_122_24), .Q(\values[1] [10]), 
      .QN());
   DFF_X1 \values_reg[1][9]  (.D(values[9]), .CK(n_122_24), .Q(\values[1] [9]), 
      .QN());
   DFF_X1 \values_reg[1][8]  (.D(values[8]), .CK(n_122_24), .Q(\values[1] [8]), 
      .QN());
   DFF_X1 \values_reg[1][7]  (.D(values[7]), .CK(n_122_24), .Q(\values[1] [7]), 
      .QN());
   DFF_X1 \values_reg[1][6]  (.D(values[6]), .CK(n_122_24), .Q(\values[1] [6]), 
      .QN());
   DFF_X1 \values_reg[1][5]  (.D(values[5]), .CK(n_122_24), .Q(\values[1] [5]), 
      .QN());
   DFF_X1 \values_reg[1][4]  (.D(values[4]), .CK(n_122_24), .Q(\values[1] [4]), 
      .QN());
   DFF_X1 \values_reg[1][3]  (.D(values[3]), .CK(n_122_24), .Q(\values[1] [3]), 
      .QN());
   DFF_X1 \values_reg[1][2]  (.D(values[2]), .CK(n_122_24), .Q(\values[1] [2]), 
      .QN());
   DFF_X1 \values_reg[1][1]  (.D(values[1]), .CK(n_122_24), .Q(\values[1] [1]), 
      .QN());
   DFF_X1 \values_reg[1][0]  (.D(values[0]), .CK(n_122_24), .Q(\values[1] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_values_reg[0]_reg  (.CK(clk), .E(n_0), .SE(1'b0), 
      .GCK(n_122_25));
   DFF_X1 \values_reg[0][15]  (.D(values[15]), .CK(n_122_25), .Q(\values[0] [15]), 
      .QN());
   DFF_X1 \values_reg[0][14]  (.D(values[14]), .CK(n_122_25), .Q(\values[0] [14]), 
      .QN());
   DFF_X1 \values_reg[0][13]  (.D(values[13]), .CK(n_122_25), .Q(\values[0] [13]), 
      .QN());
   DFF_X1 \values_reg[0][12]  (.D(values[12]), .CK(n_122_25), .Q(\values[0] [12]), 
      .QN());
   DFF_X1 \values_reg[0][11]  (.D(values[11]), .CK(n_122_25), .Q(\values[0] [11]), 
      .QN());
   DFF_X1 \values_reg[0][10]  (.D(values[10]), .CK(n_122_25), .Q(\values[0] [10]), 
      .QN());
   DFF_X1 \values_reg[0][9]  (.D(values[9]), .CK(n_122_25), .Q(\values[0] [9]), 
      .QN());
   DFF_X1 \values_reg[0][8]  (.D(values[8]), .CK(n_122_25), .Q(\values[0] [8]), 
      .QN());
   DFF_X1 \values_reg[0][7]  (.D(values[7]), .CK(n_122_25), .Q(\values[0] [7]), 
      .QN());
   DFF_X1 \values_reg[0][6]  (.D(values[6]), .CK(n_122_25), .Q(\values[0] [6]), 
      .QN());
   DFF_X1 \values_reg[0][5]  (.D(values[5]), .CK(n_122_25), .Q(\values[0] [5]), 
      .QN());
   DFF_X1 \values_reg[0][4]  (.D(values[4]), .CK(n_122_25), .Q(\values[0] [4]), 
      .QN());
   DFF_X1 \values_reg[0][3]  (.D(values[3]), .CK(n_122_25), .Q(\values[0] [3]), 
      .QN());
   DFF_X1 \values_reg[0][2]  (.D(values[2]), .CK(n_122_25), .Q(\values[0] [2]), 
      .QN());
   DFF_X1 \values_reg[0][1]  (.D(values[1]), .CK(n_122_25), .Q(\values[0] [1]), 
      .QN());
   DFF_X1 \values_reg[0][0]  (.D(values[0]), .CK(n_122_25), .Q(\values[0] [0]), 
      .QN());
   INV_X1 i_0_0_0 (.A(reset), .ZN(n_0_0_0));
   AND2_X1 i_0_0_1 (.A1(n_0_0_0), .A2(load_value[0]), .ZN(values[0]));
   AND2_X1 i_0_0_2 (.A1(n_0_0_0), .A2(load_value[1]), .ZN(values[1]));
   AND2_X1 i_0_0_3 (.A1(n_0_0_0), .A2(load_value[2]), .ZN(values[2]));
   AND2_X1 i_0_0_4 (.A1(n_0_0_0), .A2(load_value[3]), .ZN(values[3]));
   AND2_X1 i_0_0_5 (.A1(n_0_0_0), .A2(load_value[4]), .ZN(values[4]));
   AND2_X1 i_0_0_6 (.A1(n_0_0_0), .A2(load_value[5]), .ZN(values[5]));
   AND2_X1 i_0_0_7 (.A1(n_0_0_0), .A2(load_value[6]), .ZN(values[6]));
   AND2_X1 i_0_0_8 (.A1(n_0_0_0), .A2(load_value[7]), .ZN(values[7]));
   AND2_X1 i_0_0_9 (.A1(n_0_0_0), .A2(load_value[8]), .ZN(values[8]));
   AND2_X1 i_0_0_10 (.A1(n_0_0_0), .A2(load_value[9]), .ZN(values[9]));
   AND2_X1 i_0_0_11 (.A1(n_0_0_0), .A2(load_value[10]), .ZN(values[10]));
   AND2_X1 i_0_0_12 (.A1(n_0_0_0), .A2(load_value[11]), .ZN(values[11]));
   AND2_X1 i_0_0_13 (.A1(n_0_0_0), .A2(load_value[12]), .ZN(values[12]));
   AND2_X1 i_0_0_14 (.A1(n_0_0_0), .A2(load_value[13]), .ZN(values[13]));
   AND2_X1 i_0_0_15 (.A1(n_0_0_0), .A2(load_value[14]), .ZN(values[14]));
   AND2_X1 i_0_0_16 (.A1(n_0_0_0), .A2(load_value[15]), .ZN(values[15]));
   NOR4_X1 i_0_0_17 (.A1(load_address[14]), .A2(load_address[13]), .A3(
      load_address[12]), .A4(load_address[11]), .ZN(n_0_0_1));
   NOR4_X1 i_0_0_18 (.A1(load_address[10]), .A2(load_address[9]), .A3(
      load_address[8]), .A4(load_address[7]), .ZN(n_0_0_2));
   INV_X1 i_0_0_19 (.A(load_address[15]), .ZN(n_0_0_3));
   AND4_X1 i_0_0_20 (.A1(n_0_0_1), .A2(n_0_0_2), .A3(n_0_0_3), .A4(load_en), 
      .ZN(n_0_0_4));
   INV_X1 i_0_0_21 (.A(load_address[1]), .ZN(n_0_0_5));
   NAND2_X1 i_0_0_22 (.A1(n_0_0_4), .A2(n_0_0_5), .ZN(n_0_0_6));
   NOR2_X1 i_0_0_23 (.A1(n_0_0_6), .A2(load_address[3]), .ZN(n_0_0_7));
   NOR2_X1 i_0_0_24 (.A1(load_address[6]), .A2(load_address[5]), .ZN(n_0_0_8));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_7), .A2(n_0_0_8), .ZN(n_0_0_9));
   INV_X1 i_0_0_26 (.A(load_address[4]), .ZN(n_0_0_10));
   INV_X1 i_0_0_27 (.A(load_address[2]), .ZN(n_0_0_11));
   INV_X1 i_0_0_28 (.A(load_address[0]), .ZN(n_0_0_12));
   NAND3_X1 i_0_0_29 (.A1(n_0_0_10), .A2(n_0_0_11), .A3(n_0_0_12), .ZN(n_0_0_13));
   OAI21_X1 i_0_0_30 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_13), .ZN(n_0));
   NAND3_X1 i_0_0_31 (.A1(n_0_0_10), .A2(n_0_0_11), .A3(load_address[0]), 
      .ZN(n_0_0_14));
   OAI21_X1 i_0_0_32 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_14), .ZN(n_1));
   NAND2_X1 i_0_0_33 (.A1(n_0_0_4), .A2(load_address[1]), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_15), .A2(load_address[3]), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_16), .A2(n_0_0_8), .ZN(n_0_0_17));
   OAI21_X1 i_0_0_36 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_13), .ZN(n_2));
   OAI21_X1 i_0_0_37 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_14), .ZN(n_3));
   NAND3_X1 i_0_0_38 (.A1(n_0_0_10), .A2(n_0_0_12), .A3(load_address[2]), 
      .ZN(n_0_0_18));
   OAI21_X1 i_0_0_39 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_18), .ZN(n_4));
   NAND3_X1 i_0_0_40 (.A1(n_0_0_10), .A2(load_address[2]), .A3(load_address[0]), 
      .ZN(n_0_0_19));
   OAI21_X1 i_0_0_41 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_19), .ZN(n_5));
   OAI21_X1 i_0_0_42 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_18), .ZN(n_6));
   OAI21_X1 i_0_0_43 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_19), .ZN(n_7));
   INV_X1 i_0_0_44 (.A(load_address[3]), .ZN(n_0_0_20));
   NOR2_X1 i_0_0_45 (.A1(n_0_0_6), .A2(n_0_0_20), .ZN(n_0_0_21));
   NAND2_X1 i_0_0_46 (.A1(n_0_0_21), .A2(n_0_0_8), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_47 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_13), .ZN(n_8));
   OAI21_X1 i_0_0_48 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_14), .ZN(n_9));
   NOR2_X1 i_0_0_49 (.A1(n_0_0_15), .A2(n_0_0_20), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_23), .A2(n_0_0_8), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_51 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_13), .ZN(n_10));
   OAI21_X1 i_0_0_52 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_14), .ZN(n_11));
   OAI21_X1 i_0_0_53 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_18), .ZN(n_12));
   OAI21_X1 i_0_0_54 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_19), .ZN(n_13));
   OAI21_X1 i_0_0_55 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_18), .ZN(n_14));
   OAI21_X1 i_0_0_56 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_19), .ZN(n_15));
   NAND3_X1 i_0_0_57 (.A1(n_0_0_12), .A2(n_0_0_11), .A3(load_address[4]), 
      .ZN(n_0_0_25));
   OAI21_X1 i_0_0_58 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_25), .ZN(n_16));
   NAND3_X1 i_0_0_59 (.A1(n_0_0_11), .A2(load_address[4]), .A3(load_address[0]), 
      .ZN(n_0_0_26));
   OAI21_X1 i_0_0_60 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_26), .ZN(n_17));
   OAI21_X1 i_0_0_61 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_25), .ZN(n_18));
   OAI21_X1 i_0_0_62 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_26), .ZN(n_19));
   NAND3_X1 i_0_0_63 (.A1(n_0_0_12), .A2(load_address[4]), .A3(load_address[2]), 
      .ZN(n_0_0_27));
   OAI21_X1 i_0_0_64 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_27), .ZN(n_20));
   NAND3_X1 i_0_0_65 (.A1(load_address[4]), .A2(load_address[2]), .A3(
      load_address[0]), .ZN(n_0_0_28));
   OAI21_X1 i_0_0_66 (.A(n_0_0_0), .B1(n_0_0_9), .B2(n_0_0_28), .ZN(n_21));
   OAI21_X1 i_0_0_67 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_27), .ZN(n_22));
   OAI21_X1 i_0_0_68 (.A(n_0_0_0), .B1(n_0_0_17), .B2(n_0_0_28), .ZN(n_23));
   OAI21_X1 i_0_0_69 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_25), .ZN(n_24));
   OAI21_X1 i_0_0_70 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_26), .ZN(n_25));
   OAI21_X1 i_0_0_71 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_25), .ZN(n_26));
   OAI21_X1 i_0_0_72 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_26), .ZN(n_27));
   OAI21_X1 i_0_0_73 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_27), .ZN(n_28));
   OAI21_X1 i_0_0_74 (.A(n_0_0_0), .B1(n_0_0_22), .B2(n_0_0_28), .ZN(n_29));
   OAI21_X1 i_0_0_75 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_27), .ZN(n_30));
   OAI21_X1 i_0_0_76 (.A(n_0_0_0), .B1(n_0_0_24), .B2(n_0_0_28), .ZN(n_31));
   INV_X1 i_0_0_77 (.A(load_address[5]), .ZN(n_0_0_29));
   NOR2_X1 i_0_0_78 (.A1(n_0_0_29), .A2(load_address[6]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_79 (.A1(n_0_0_7), .A2(n_0_0_30), .ZN(n_0_0_31));
   OAI21_X1 i_0_0_80 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_13), .ZN(n_32));
   OAI21_X1 i_0_0_81 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_14), .ZN(n_33));
   NAND2_X1 i_0_0_82 (.A1(n_0_0_16), .A2(n_0_0_30), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_83 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_13), .ZN(n_34));
   OAI21_X1 i_0_0_84 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_14), .ZN(n_35));
   OAI21_X1 i_0_0_85 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_18), .ZN(n_36));
   OAI21_X1 i_0_0_86 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_19), .ZN(n_37));
   OAI21_X1 i_0_0_87 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_18), .ZN(n_38));
   OAI21_X1 i_0_0_88 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_19), .ZN(n_39));
   NAND2_X1 i_0_0_89 (.A1(n_0_0_21), .A2(n_0_0_30), .ZN(n_0_0_33));
   OAI21_X1 i_0_0_90 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_13), .ZN(n_40));
   OAI21_X1 i_0_0_91 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_14), .ZN(n_41));
   NAND2_X1 i_0_0_92 (.A1(n_0_0_23), .A2(n_0_0_30), .ZN(n_0_0_34));
   OAI21_X1 i_0_0_93 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_13), .ZN(n_42));
   OAI21_X1 i_0_0_94 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_14), .ZN(n_43));
   OAI21_X1 i_0_0_95 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_18), .ZN(n_44));
   OAI21_X1 i_0_0_96 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_19), .ZN(n_45));
   OAI21_X1 i_0_0_97 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_18), .ZN(n_46));
   OAI21_X1 i_0_0_98 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_19), .ZN(n_47));
   OAI21_X1 i_0_0_99 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_25), .ZN(n_48));
   OAI21_X1 i_0_0_100 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_26), .ZN(n_49));
   OAI21_X1 i_0_0_101 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_25), .ZN(n_50));
   OAI21_X1 i_0_0_102 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_26), .ZN(n_51));
   OAI21_X1 i_0_0_103 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_27), .ZN(n_52));
   OAI21_X1 i_0_0_104 (.A(n_0_0_0), .B1(n_0_0_31), .B2(n_0_0_28), .ZN(n_53));
   OAI21_X1 i_0_0_105 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_27), .ZN(n_54));
   OAI21_X1 i_0_0_106 (.A(n_0_0_0), .B1(n_0_0_32), .B2(n_0_0_28), .ZN(n_55));
   OAI21_X1 i_0_0_107 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_25), .ZN(n_56));
   OAI21_X1 i_0_0_108 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_26), .ZN(n_57));
   OAI21_X1 i_0_0_109 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_25), .ZN(n_58));
   OAI21_X1 i_0_0_110 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_26), .ZN(n_59));
   OAI21_X1 i_0_0_111 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_27), .ZN(n_60));
   OAI21_X1 i_0_0_112 (.A(n_0_0_0), .B1(n_0_0_33), .B2(n_0_0_28), .ZN(n_61));
   OAI21_X1 i_0_0_113 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_27), .ZN(n_62));
   OAI21_X1 i_0_0_114 (.A(n_0_0_0), .B1(n_0_0_34), .B2(n_0_0_28), .ZN(n_63));
   INV_X1 i_0_0_115 (.A(load_address[6]), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_116 (.A1(n_0_0_35), .A2(load_address[5]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_117 (.A1(n_0_0_7), .A2(n_0_0_36), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_118 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_13), .ZN(n_64));
   OAI21_X1 i_0_0_119 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_14), .ZN(n_65));
   NAND2_X1 i_0_0_120 (.A1(n_0_0_16), .A2(n_0_0_36), .ZN(n_0_0_38));
   OAI21_X1 i_0_0_121 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_13), .ZN(n_66));
   OAI21_X1 i_0_0_122 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_14), .ZN(n_67));
   OAI21_X1 i_0_0_123 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_18), .ZN(n_68));
   OAI21_X1 i_0_0_124 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_19), .ZN(n_69));
   OAI21_X1 i_0_0_125 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_18), .ZN(n_70));
   OAI21_X1 i_0_0_126 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_19), .ZN(n_71));
   NAND2_X1 i_0_0_127 (.A1(n_0_0_21), .A2(n_0_0_36), .ZN(n_0_0_39));
   OAI21_X1 i_0_0_128 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_13), .ZN(n_72));
   OAI21_X1 i_0_0_129 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_14), .ZN(n_73));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_23), .A2(n_0_0_36), .ZN(n_0_0_40));
   OAI21_X1 i_0_0_131 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_13), .ZN(n_74));
   OAI21_X1 i_0_0_132 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_14), .ZN(n_75));
   OAI21_X1 i_0_0_133 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_18), .ZN(n_76));
   OAI21_X1 i_0_0_134 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_19), .ZN(n_77));
   OAI21_X1 i_0_0_135 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_18), .ZN(n_78));
   OAI21_X1 i_0_0_136 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_19), .ZN(n_79));
   OAI21_X1 i_0_0_137 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_25), .ZN(n_80));
   OAI21_X1 i_0_0_138 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_26), .ZN(n_81));
   OAI21_X1 i_0_0_139 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_25), .ZN(n_82));
   OAI21_X1 i_0_0_140 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_26), .ZN(n_83));
   OAI21_X1 i_0_0_141 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_27), .ZN(n_84));
   OAI21_X1 i_0_0_142 (.A(n_0_0_0), .B1(n_0_0_37), .B2(n_0_0_28), .ZN(n_85));
   OAI21_X1 i_0_0_143 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_27), .ZN(n_86));
   OAI21_X1 i_0_0_144 (.A(n_0_0_0), .B1(n_0_0_38), .B2(n_0_0_28), .ZN(n_87));
   OAI21_X1 i_0_0_145 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_25), .ZN(n_88));
   OAI21_X1 i_0_0_146 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_26), .ZN(n_89));
   OAI21_X1 i_0_0_147 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_25), .ZN(n_90));
   OAI21_X1 i_0_0_148 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_26), .ZN(n_91));
   OAI21_X1 i_0_0_149 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_27), .ZN(n_92));
   OAI21_X1 i_0_0_150 (.A(n_0_0_0), .B1(n_0_0_39), .B2(n_0_0_28), .ZN(n_93));
   OAI21_X1 i_0_0_151 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_27), .ZN(n_94));
   OAI21_X1 i_0_0_152 (.A(n_0_0_0), .B1(n_0_0_40), .B2(n_0_0_28), .ZN(n_95));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_35), .A2(n_0_0_29), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_154 (.A1(n_0_0_7), .A2(n_0_0_41), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_155 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_13), .ZN(n_96));
   OAI21_X1 i_0_0_156 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_14), .ZN(n_97));
   NAND2_X1 i_0_0_157 (.A1(n_0_0_16), .A2(n_0_0_41), .ZN(n_0_0_43));
   OAI21_X1 i_0_0_158 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_13), .ZN(n_98));
   OAI21_X1 i_0_0_159 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_14), .ZN(n_99));
   OAI21_X1 i_0_0_160 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_18), .ZN(n_100));
   OAI21_X1 i_0_0_161 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_19), .ZN(n_101));
   OAI21_X1 i_0_0_162 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_18), .ZN(n_102));
   OAI21_X1 i_0_0_163 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_19), .ZN(n_103));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_21), .A2(n_0_0_41), .ZN(n_0_0_44));
   OAI21_X1 i_0_0_165 (.A(n_0_0_0), .B1(n_0_0_44), .B2(n_0_0_13), .ZN(n_104));
   OAI21_X1 i_0_0_166 (.A(n_0_0_0), .B1(n_0_0_44), .B2(n_0_0_14), .ZN(n_105));
   NAND2_X1 i_0_0_167 (.A1(n_0_0_23), .A2(n_0_0_41), .ZN(n_0_0_45));
   OAI21_X1 i_0_0_168 (.A(n_0_0_0), .B1(n_0_0_45), .B2(n_0_0_13), .ZN(n_106));
   OAI21_X1 i_0_0_169 (.A(n_0_0_0), .B1(n_0_0_45), .B2(n_0_0_14), .ZN(n_107));
   OAI21_X1 i_0_0_170 (.A(n_0_0_0), .B1(n_0_0_44), .B2(n_0_0_18), .ZN(n_108));
   OAI21_X1 i_0_0_171 (.A(n_0_0_0), .B1(n_0_0_44), .B2(n_0_0_19), .ZN(n_109));
   OAI21_X1 i_0_0_172 (.A(n_0_0_0), .B1(n_0_0_45), .B2(n_0_0_18), .ZN(n_110));
   OAI21_X1 i_0_0_173 (.A(n_0_0_0), .B1(n_0_0_45), .B2(n_0_0_19), .ZN(n_111));
   OAI21_X1 i_0_0_174 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_25), .ZN(n_112));
   OAI21_X1 i_0_0_175 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_26), .ZN(n_113));
   OAI21_X1 i_0_0_176 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_25), .ZN(n_114));
   OAI21_X1 i_0_0_177 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_26), .ZN(n_115));
   OAI21_X1 i_0_0_178 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_27), .ZN(n_116));
   OAI21_X1 i_0_0_179 (.A(n_0_0_0), .B1(n_0_0_42), .B2(n_0_0_28), .ZN(n_117));
   OAI21_X1 i_0_0_180 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_27), .ZN(n_118));
   OAI21_X1 i_0_0_181 (.A(n_0_0_0), .B1(n_0_0_43), .B2(n_0_0_28), .ZN(n_119));
endmodule
