
// 	Wed May  5 23:39:23 2021
//	vlsi
//	localhost.localdomain

module Neuron_Layer (clk, load_en, load_value, load_address, reset, \o_values[0] , 
    \o_values[1] , \o_values[2] , \o_values[3] , \o_values[4] , \o_values[5] , \o_values[6] , 
    \o_values[7] , \o_values[8] , \o_values[9] , \o_values[10] , \o_values[11] , 
    \o_values[12] , \o_values[13] , \o_values[14] , \o_values[15] , \o_values[16] , 
    \o_values[17] , \o_values[18] , \o_values[19] , \o_values[20] , \o_values[21] , 
    \o_values[22] , \o_values[23] , \o_values[24] , \o_values[25] , \o_values[26] , 
    \o_values[27] , \o_values[28] , \o_values[29] , \o_values[30] , \o_values[31] , 
    \o_values[32] , \o_values[33] , \o_values[34] , \o_values[35] , \o_values[36] , 
    \o_values[37] , \o_values[38] , \o_values[39] , \o_values[40] , \o_values[41] , 
    \o_values[42] , \o_values[43] , \o_values[44] , \o_values[45] , \o_values[46] , 
    \o_values[47] , \o_values[48] , \o_values[49] , \o_values[50] , \o_values[51] , 
    \o_values[52] , \o_values[53] , \o_values[54] , \o_values[55] , \o_values[56] , 
    \o_values[57] , \o_values[58] , \o_values[59] , \o_values[60] , \o_values[61] , 
    \o_values[62] , \o_values[63] , \o_values[64] , \o_values[65] , \o_values[66] , 
    \o_values[67] , \o_values[68] , \o_values[69] , \o_values[70] , \o_values[71] , 
    \o_values[72] , \o_values[73] , \o_values[74] , \o_values[75] , \o_values[76] , 
    \o_values[77] , \o_values[78] , \o_values[79] , \o_values[80] , \o_values[81] , 
    \o_values[82] , \o_values[83] );

output [15:0] \o_values[0] ;
output [15:0] \o_values[10] ;
output [15:0] \o_values[11] ;
output [15:0] \o_values[12] ;
output [15:0] \o_values[13] ;
output [15:0] \o_values[14] ;
output [15:0] \o_values[15] ;
output [15:0] \o_values[16] ;
output [15:0] \o_values[17] ;
output [15:0] \o_values[18] ;
output [15:0] \o_values[19] ;
output [15:0] \o_values[1] ;
output [15:0] \o_values[20] ;
output [15:0] \o_values[21] ;
output [15:0] \o_values[22] ;
output [15:0] \o_values[23] ;
output [15:0] \o_values[24] ;
output [15:0] \o_values[25] ;
output [15:0] \o_values[26] ;
output [15:0] \o_values[27] ;
output [15:0] \o_values[28] ;
output [15:0] \o_values[29] ;
output [15:0] \o_values[2] ;
output [15:0] \o_values[30] ;
output [15:0] \o_values[31] ;
output [15:0] \o_values[32] ;
output [15:0] \o_values[33] ;
output [15:0] \o_values[34] ;
output [15:0] \o_values[35] ;
output [15:0] \o_values[36] ;
output [15:0] \o_values[37] ;
output [15:0] \o_values[38] ;
output [15:0] \o_values[39] ;
output [15:0] \o_values[3] ;
output [15:0] \o_values[40] ;
output [15:0] \o_values[41] ;
output [15:0] \o_values[42] ;
output [15:0] \o_values[43] ;
output [15:0] \o_values[44] ;
output [15:0] \o_values[45] ;
output [15:0] \o_values[46] ;
output [15:0] \o_values[47] ;
output [15:0] \o_values[48] ;
output [15:0] \o_values[49] ;
output [15:0] \o_values[4] ;
output [15:0] \o_values[50] ;
output [15:0] \o_values[51] ;
output [15:0] \o_values[52] ;
output [15:0] \o_values[53] ;
output [15:0] \o_values[54] ;
output [15:0] \o_values[55] ;
output [15:0] \o_values[56] ;
output [15:0] \o_values[57] ;
output [15:0] \o_values[58] ;
output [15:0] \o_values[59] ;
output [15:0] \o_values[5] ;
output [15:0] \o_values[60] ;
output [15:0] \o_values[61] ;
output [15:0] \o_values[62] ;
output [15:0] \o_values[63] ;
output [15:0] \o_values[64] ;
output [15:0] \o_values[65] ;
output [15:0] \o_values[66] ;
output [15:0] \o_values[67] ;
output [15:0] \o_values[68] ;
output [15:0] \o_values[69] ;
output [15:0] \o_values[6] ;
output [15:0] \o_values[70] ;
output [15:0] \o_values[71] ;
output [15:0] \o_values[72] ;
output [15:0] \o_values[73] ;
output [15:0] \o_values[74] ;
output [15:0] \o_values[75] ;
output [15:0] \o_values[76] ;
output [15:0] \o_values[77] ;
output [15:0] \o_values[78] ;
output [15:0] \o_values[79] ;
output [15:0] \o_values[7] ;
output [15:0] \o_values[80] ;
output [15:0] \o_values[81] ;
output [15:0] \o_values[82] ;
output [15:0] \o_values[83] ;
output [15:0] \o_values[8] ;
output [15:0] \o_values[9] ;
input clk;
input [15:0] load_address;
input load_en;
input [15:0] load_value;
input reset;
wire n_0_84;
wire n_0_85;
wire n_0_86;
wire n_0_87;
wire n_0_88;
wire n_0_89;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_93;
wire n_0_94;
wire n_0_95;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_103;
wire n_0_104;
wire n_0_105;
wire n_0_106;
wire n_0_107;
wire n_0_108;
wire n_0_109;
wire n_0_110;
wire n_0_111;
wire n_0_112;
wire n_0_113;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_139;
wire n_0_140;
wire n_0_141;
wire n_0_142;
wire n_0_143;
wire n_0_144;
wire n_0_145;
wire n_0_146;
wire n_0_147;
wire n_0_148;
wire n_0_149;
wire n_0_150;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire \t_o_values[14] ;
wire \t_o_values[15] ;
wire \t_o_values[13] ;
wire \t_o_values[12] ;
wire \t_o_values[11] ;
wire \t_o_values[10] ;
wire \t_o_values[9] ;
wire \t_o_values[8] ;
wire \t_o_values[7] ;
wire \t_o_values[6] ;
wire \t_o_values[5] ;
wire \t_o_values[4] ;
wire \t_o_values[3] ;
wire \t_o_values[2] ;
wire \t_o_values[1] ;
wire \t_o_values[0] ;
wire n_0_83;
wire n_0_82;
wire n_0_81;
wire n_0_80;
wire n_0_0_0;
wire n_0_79;
wire n_0_78;
wire n_0_77;
wire n_0_76;
wire n_0_0_1;
wire n_0_75;
wire n_0_74;
wire n_0_73;
wire n_0_72;
wire n_0_0_2;
wire n_0_71;
wire n_0_70;
wire n_0_69;
wire n_0_68;
wire n_0_0_3;
wire n_0_67;
wire n_0_66;
wire n_0_65;
wire n_0_64;
wire n_0_63;
wire n_0_62;
wire n_0_61;
wire n_0_60;
wire n_0_0_4;
wire n_0_59;
wire n_0_58;
wire n_0_57;
wire n_0_56;
wire n_0_0_5;
wire n_0_55;
wire n_0_54;
wire n_0_53;
wire n_0_52;
wire n_0_0_6;
wire n_0_51;
wire n_0_50;
wire n_0_49;
wire n_0_48;
wire n_0_0_7;
wire n_0_47;
wire n_0_46;
wire n_0_45;
wire n_0_44;
wire n_0_0_8;
wire n_0_43;
wire n_0_42;
wire n_0_41;
wire n_0_40;
wire n_0_0_9;
wire n_0_39;
wire n_0_38;
wire n_0_37;
wire n_0_36;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_35;
wire n_0_34;
wire n_0_33;
wire n_0_32;
wire n_0_0_12;
wire n_0_31;
wire n_0_30;
wire n_0_29;
wire n_0_28;
wire n_0_0_13;
wire n_0_27;
wire n_0_26;
wire n_0_25;
wire n_0_24;
wire n_0_0_14;
wire n_0_23;
wire n_0_0_15;
wire n_0_22;
wire n_0_0_16;
wire n_0_21;
wire n_0_0_17;
wire n_0_20;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_19;
wire n_0_18;
wire n_0_17;
wire n_0_16;
wire n_0_15;
wire n_0_14;
wire n_0_13;
wire n_0_12;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_11;
wire n_0_10;
wire n_0_9;
wire n_0_8;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_7;
wire n_0_0_25;
wire n_0_6;
wire n_0_0_26;
wire n_0_5;
wire n_0_0_27;
wire n_0_4;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_3;
wire n_0_0_33;
wire n_0_2;
wire n_0_0_34;
wire n_0_1;
wire n_0_0_35;
wire n_0_0;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire sps__n1;
wire sps__n4;
wire sps__n7;
wire sps__n10;
wire sps__n13;
wire sps__n16;
wire sps__n19;
wire sps__n22;
wire sps__n25;
wire sps__n28;
wire sps__n31;
wire sps__n34;
wire sps__n37;


INV_X4 i_0_0_152 (.ZN (n_0_0_52), .A (reset));
INV_X1 i_0_0_151 (.ZN (n_0_0_51), .A (load_en));
INV_X1 i_0_0_150 (.ZN (n_0_0_50), .A (load_address[4]));
INV_X1 i_0_0_149 (.ZN (n_0_0_49), .A (load_address[3]));
INV_X1 i_0_0_148 (.ZN (n_0_0_48), .A (load_address[2]));
INV_X1 i_0_0_147 (.ZN (n_0_0_47), .A (load_address[1]));
INV_X1 i_0_0_146 (.ZN (n_0_0_46), .A (load_address[0]));
NAND2_X1 i_0_0_145 (.ZN (n_0_0_45), .A1 (load_address[1]), .A2 (load_address[0]));
OR4_X1 i_0_0_144 (.ZN (n_0_0_44), .A1 (n_0_0_51), .A2 (load_address[15]), .A3 (load_address[14]), .A4 (load_address[13]));
OR4_X1 i_0_0_143 (.ZN (n_0_0_43), .A1 (load_address[12]), .A2 (load_address[11]), .A3 (load_address[10]), .A4 (load_address[9]));
NOR2_X1 i_0_0_142 (.ZN (n_0_0_42), .A1 (load_address[3]), .A2 (load_address[2]));
NAND2_X1 i_0_0_141 (.ZN (n_0_0_41), .A1 (n_0_0_49), .A2 (n_0_0_48));
NOR2_X1 i_0_0_140 (.ZN (n_0_0_40), .A1 (n_0_0_50), .A2 (load_address[5]));
NAND2_X1 i_0_0_139 (.ZN (n_0_0_39), .A1 (n_0_0_42), .A2 (n_0_0_40));
NOR4_X1 i_0_0_138 (.ZN (n_0_0_38), .A1 (n_0_0_44), .A2 (n_0_0_43), .A3 (load_address[8]), .A4 (load_address[7]));
INV_X1 i_0_0_137 (.ZN (n_0_0_37), .A (n_0_0_38));
NAND4_X1 i_0_0_136 (.ZN (n_0_0_36), .A1 (load_address[6]), .A2 (n_0_0_42), .A3 (n_0_0_40), .A4 (n_0_0_38));
OAI21_X1 i_0_0_135 (.ZN (n_0_0), .A (n_0_0_52), .B1 (n_0_0_45), .B2 (n_0_0_36));
NAND2_X1 i_0_0_134 (.ZN (n_0_0_35), .A1 (n_0_0_46), .A2 (load_address[1]));
OAI21_X1 i_0_0_133 (.ZN (n_0_1), .A (n_0_0_52), .B1 (n_0_0_36), .B2 (n_0_0_35));
NAND2_X1 i_0_0_132 (.ZN (n_0_0_34), .A1 (n_0_0_47), .A2 (load_address[0]));
OAI21_X1 i_0_0_131 (.ZN (n_0_2), .A (n_0_0_52), .B1 (n_0_0_36), .B2 (n_0_0_34));
NAND2_X1 i_0_0_130 (.ZN (n_0_0_33), .A1 (n_0_0_47), .A2 (n_0_0_46));
OAI21_X1 i_0_0_129 (.ZN (n_0_3), .A (n_0_0_52), .B1 (n_0_0_36), .B2 (n_0_0_33));
NOR2_X1 i_0_0_128 (.ZN (n_0_0_32), .A1 (n_0_0_49), .A2 (n_0_0_48));
NAND2_X1 i_0_0_127 (.ZN (n_0_0_31), .A1 (load_address[3]), .A2 (load_address[2]));
NOR2_X1 i_0_0_126 (.ZN (n_0_0_30), .A1 (load_address[5]), .A2 (load_address[4]));
NAND3_X1 i_0_0_125 (.ZN (n_0_0_29), .A1 (load_address[6]), .A2 (n_0_0_38), .A3 (n_0_0_30));
OR2_X1 i_0_0_124 (.ZN (n_0_0_28), .A1 (n_0_0_45), .A2 (n_0_0_29));
OAI21_X1 i_0_0_123 (.ZN (n_0_4), .A (n_0_0_52), .B1 (n_0_0_31), .B2 (n_0_0_28));
OR2_X1 i_0_0_122 (.ZN (n_0_0_27), .A1 (n_0_0_35), .A2 (n_0_0_29));
OAI21_X1 i_0_0_121 (.ZN (n_0_5), .A (n_0_0_52), .B1 (n_0_0_31), .B2 (n_0_0_27));
OR2_X1 i_0_0_120 (.ZN (n_0_0_26), .A1 (n_0_0_34), .A2 (n_0_0_29));
OAI21_X1 i_0_0_119 (.ZN (n_0_6), .A (n_0_0_52), .B1 (n_0_0_31), .B2 (n_0_0_26));
OR2_X1 i_0_0_118 (.ZN (n_0_0_25), .A1 (n_0_0_33), .A2 (n_0_0_29));
OAI21_X1 i_0_0_117 (.ZN (n_0_7), .A (n_0_0_52), .B1 (n_0_0_31), .B2 (n_0_0_25));
NOR2_X1 i_0_0_116 (.ZN (n_0_0_24), .A1 (n_0_0_49), .A2 (load_address[2]));
NAND2_X1 i_0_0_115 (.ZN (n_0_0_23), .A1 (n_0_0_48), .A2 (load_address[3]));
OAI21_X1 i_0_0_114 (.ZN (n_0_8), .A (n_0_0_52), .B1 (n_0_0_28), .B2 (n_0_0_23));
OAI21_X1 i_0_0_113 (.ZN (n_0_9), .A (n_0_0_52), .B1 (n_0_0_27), .B2 (n_0_0_23));
OAI21_X1 i_0_0_112 (.ZN (n_0_10), .A (n_0_0_52), .B1 (n_0_0_26), .B2 (n_0_0_23));
OAI21_X1 i_0_0_111 (.ZN (n_0_11), .A (n_0_0_52), .B1 (n_0_0_25), .B2 (n_0_0_23));
NOR2_X1 i_0_0_110 (.ZN (n_0_0_22), .A1 (n_0_0_48), .A2 (load_address[3]));
NAND2_X1 i_0_0_109 (.ZN (n_0_0_21), .A1 (n_0_0_49), .A2 (load_address[2]));
OAI21_X1 i_0_0_108 (.ZN (n_0_12), .A (n_0_0_52), .B1 (n_0_0_28), .B2 (n_0_0_21));
OAI21_X1 i_0_0_107 (.ZN (n_0_13), .A (n_0_0_52), .B1 (n_0_0_27), .B2 (n_0_0_21));
OAI21_X1 i_0_0_106 (.ZN (n_0_14), .A (n_0_0_52), .B1 (n_0_0_26), .B2 (n_0_0_21));
OAI21_X1 i_0_0_105 (.ZN (n_0_15), .A (n_0_0_52), .B1 (n_0_0_25), .B2 (n_0_0_21));
OAI21_X1 i_0_0_104 (.ZN (n_0_16), .A (n_0_0_52), .B1 (n_0_0_41), .B2 (n_0_0_28));
OAI21_X1 i_0_0_103 (.ZN (n_0_17), .A (n_0_0_52), .B1 (n_0_0_41), .B2 (n_0_0_27));
OAI21_X1 i_0_0_102 (.ZN (n_0_18), .A (n_0_0_52), .B1 (n_0_0_41), .B2 (n_0_0_26));
OAI21_X1 i_0_0_101 (.ZN (n_0_19), .A (n_0_0_52), .B1 (n_0_0_41), .B2 (n_0_0_25));
NAND3_X1 i_0_0_100 (.ZN (n_0_0_20), .A1 (load_address[5]), .A2 (load_address[4]), .A3 (n_0_0_32));
NOR2_X1 i_0_0_99 (.ZN (n_0_0_19), .A1 (n_0_0_37), .A2 (load_address[6]));
NAND3_X1 i_0_0_98 (.ZN (n_0_0_18), .A1 (load_address[1]), .A2 (load_address[0]), .A3 (n_0_0_19));
OAI21_X1 i_0_0_97 (.ZN (n_0_20), .A (n_0_0_52), .B1 (n_0_0_20), .B2 (n_0_0_18));
NAND3_X1 i_0_0_96 (.ZN (n_0_0_17), .A1 (load_address[1]), .A2 (n_0_0_19), .A3 (n_0_0_46));
OAI21_X1 i_0_0_95 (.ZN (n_0_21), .A (n_0_0_52), .B1 (n_0_0_20), .B2 (n_0_0_17));
NAND3_X1 i_0_0_94 (.ZN (n_0_0_16), .A1 (n_0_0_19), .A2 (n_0_0_47), .A3 (load_address[0]));
OAI21_X1 i_0_0_93 (.ZN (n_0_22), .A (n_0_0_52), .B1 (n_0_0_20), .B2 (n_0_0_16));
NAND3_X1 i_0_0_92 (.ZN (n_0_0_15), .A1 (n_0_0_19), .A2 (n_0_0_46), .A3 (n_0_0_47));
OAI21_X1 i_0_0_91 (.ZN (n_0_23), .A (n_0_0_52), .B1 (n_0_0_20), .B2 (n_0_0_15));
NAND3_X1 i_0_0_90 (.ZN (n_0_0_14), .A1 (load_address[5]), .A2 (load_address[4]), .A3 (n_0_0_24));
OAI21_X1 i_0_0_89 (.ZN (n_0_24), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_14));
OAI21_X1 i_0_0_88 (.ZN (n_0_25), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_14));
OAI21_X1 i_0_0_87 (.ZN (n_0_26), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_14));
OAI21_X1 i_0_0_86 (.ZN (n_0_27), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_14));
NAND3_X1 i_0_0_85 (.ZN (n_0_0_13), .A1 (load_address[5]), .A2 (load_address[4]), .A3 (n_0_0_22));
OAI21_X1 i_0_0_84 (.ZN (n_0_28), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_13));
OAI21_X1 i_0_0_83 (.ZN (n_0_29), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_13));
OAI21_X1 i_0_0_82 (.ZN (n_0_30), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_13));
OAI21_X1 i_0_0_81 (.ZN (n_0_31), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_13));
NAND3_X1 i_0_0_80 (.ZN (n_0_0_12), .A1 (load_address[5]), .A2 (load_address[4]), .A3 (n_0_0_42));
OAI21_X1 i_0_0_79 (.ZN (n_0_32), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_12));
OAI21_X1 i_0_0_78 (.ZN (n_0_33), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_12));
OAI21_X1 i_0_0_77 (.ZN (n_0_34), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_12));
OAI21_X1 i_0_0_76 (.ZN (n_0_35), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_12));
AND2_X1 i_0_0_75 (.ZN (n_0_0_11), .A1 (n_0_0_50), .A2 (load_address[5]));
NAND2_X1 i_0_0_74 (.ZN (n_0_0_10), .A1 (n_0_0_32), .A2 (n_0_0_11));
OAI21_X1 i_0_0_73 (.ZN (n_0_36), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_10));
OAI21_X1 i_0_0_72 (.ZN (n_0_37), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_10));
OAI21_X1 i_0_0_71 (.ZN (n_0_38), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_10));
OAI21_X1 i_0_0_70 (.ZN (n_0_39), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_10));
NAND2_X1 i_0_0_69 (.ZN (n_0_0_9), .A1 (n_0_0_24), .A2 (n_0_0_11));
OAI21_X1 i_0_0_68 (.ZN (n_0_40), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_9));
OAI21_X1 i_0_0_67 (.ZN (n_0_41), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_9));
OAI21_X1 i_0_0_66 (.ZN (n_0_42), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_9));
OAI21_X1 i_0_0_65 (.ZN (n_0_43), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_9));
NAND2_X1 i_0_0_64 (.ZN (n_0_0_8), .A1 (n_0_0_22), .A2 (n_0_0_11));
OAI21_X1 i_0_0_63 (.ZN (n_0_44), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_8));
OAI21_X1 i_0_0_62 (.ZN (n_0_45), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_8));
OAI21_X1 i_0_0_61 (.ZN (n_0_46), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_8));
OAI21_X1 i_0_0_60 (.ZN (n_0_47), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_8));
NAND2_X1 i_0_0_59 (.ZN (n_0_0_7), .A1 (n_0_0_42), .A2 (n_0_0_11));
OAI21_X1 i_0_0_58 (.ZN (n_0_48), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_7));
OAI21_X1 i_0_0_57 (.ZN (n_0_49), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_7));
OAI21_X1 i_0_0_56 (.ZN (n_0_50), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_7));
OAI21_X1 i_0_0_55 (.ZN (n_0_51), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_7));
NAND2_X1 i_0_0_54 (.ZN (n_0_0_6), .A1 (n_0_0_40), .A2 (n_0_0_32));
OAI21_X1 i_0_0_53 (.ZN (n_0_52), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_6));
OAI21_X1 i_0_0_52 (.ZN (n_0_53), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_6));
OAI21_X1 i_0_0_51 (.ZN (n_0_54), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_6));
OAI21_X1 i_0_0_50 (.ZN (n_0_55), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_6));
NAND2_X1 i_0_0_49 (.ZN (n_0_0_5), .A1 (n_0_0_40), .A2 (n_0_0_24));
OAI21_X1 i_0_0_48 (.ZN (n_0_56), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_5));
OAI21_X1 i_0_0_47 (.ZN (n_0_57), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_5));
OAI21_X1 i_0_0_46 (.ZN (n_0_58), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_5));
OAI21_X1 i_0_0_45 (.ZN (n_0_59), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_5));
NAND2_X1 i_0_0_44 (.ZN (n_0_0_4), .A1 (n_0_0_40), .A2 (n_0_0_22));
OAI21_X1 i_0_0_43 (.ZN (n_0_60), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_4));
OAI21_X1 i_0_0_42 (.ZN (n_0_61), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_4));
OAI21_X1 i_0_0_41 (.ZN (n_0_62), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_4));
OAI21_X1 i_0_0_40 (.ZN (n_0_63), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_4));
OAI21_X1 i_0_0_39 (.ZN (n_0_64), .A (n_0_0_52), .B1 (n_0_0_39), .B2 (n_0_0_18));
OAI21_X1 i_0_0_38 (.ZN (n_0_65), .A (n_0_0_52), .B1 (n_0_0_39), .B2 (n_0_0_17));
OAI21_X1 i_0_0_37 (.ZN (n_0_66), .A (n_0_0_52), .B1 (n_0_0_39), .B2 (n_0_0_16));
OAI21_X1 i_0_0_36 (.ZN (n_0_67), .A (n_0_0_52), .B1 (n_0_0_39), .B2 (n_0_0_15));
NAND2_X1 i_0_0_35 (.ZN (n_0_0_3), .A1 (n_0_0_32), .A2 (n_0_0_30));
OAI21_X1 i_0_0_34 (.ZN (n_0_68), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_3));
OAI21_X1 i_0_0_33 (.ZN (n_0_69), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_3));
OAI21_X1 i_0_0_32 (.ZN (n_0_70), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_3));
OAI21_X1 i_0_0_31 (.ZN (n_0_71), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_3));
NAND2_X1 i_0_0_30 (.ZN (n_0_0_2), .A1 (n_0_0_30), .A2 (n_0_0_24));
OAI21_X1 i_0_0_29 (.ZN (n_0_72), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_2));
OAI21_X1 i_0_0_28 (.ZN (n_0_73), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_2));
OAI21_X1 i_0_0_27 (.ZN (n_0_74), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_2));
OAI21_X1 i_0_0_26 (.ZN (n_0_75), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_2));
NAND2_X1 i_0_0_25 (.ZN (n_0_0_1), .A1 (n_0_0_30), .A2 (n_0_0_22));
OAI21_X1 i_0_0_24 (.ZN (n_0_76), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_1));
OAI21_X1 i_0_0_23 (.ZN (n_0_77), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_1));
OAI21_X1 i_0_0_22 (.ZN (n_0_78), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_1));
OAI21_X1 i_0_0_21 (.ZN (n_0_79), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_1));
NAND2_X1 i_0_0_20 (.ZN (n_0_0_0), .A1 (n_0_0_42), .A2 (n_0_0_30));
OAI21_X1 i_0_0_19 (.ZN (n_0_80), .A (n_0_0_52), .B1 (n_0_0_18), .B2 (n_0_0_0));
OAI21_X1 i_0_0_18 (.ZN (n_0_81), .A (n_0_0_52), .B1 (n_0_0_17), .B2 (n_0_0_0));
OAI21_X1 i_0_0_17 (.ZN (n_0_82), .A (n_0_0_52), .B1 (n_0_0_16), .B2 (n_0_0_0));
OAI21_X1 i_0_0_16 (.ZN (n_0_83), .A (n_0_0_52), .B1 (n_0_0_15), .B2 (n_0_0_0));
AND2_X1 i_0_0_15 (.ZN (\t_o_values[15] ), .A1 (n_0_0_52), .A2 (load_value[15]));
AND2_X1 i_0_0_14 (.ZN (\t_o_values[14] ), .A1 (n_0_0_52), .A2 (load_value[14]));
AND2_X1 i_0_0_13 (.ZN (\t_o_values[13] ), .A1 (n_0_0_52), .A2 (load_value[13]));
AND2_X1 i_0_0_12 (.ZN (\t_o_values[12] ), .A1 (n_0_0_52), .A2 (load_value[12]));
AND2_X1 i_0_0_11 (.ZN (\t_o_values[11] ), .A1 (n_0_0_52), .A2 (load_value[11]));
AND2_X1 i_0_0_10 (.ZN (\t_o_values[10] ), .A1 (n_0_0_52), .A2 (load_value[10]));
AND2_X1 i_0_0_9 (.ZN (\t_o_values[9] ), .A1 (n_0_0_52), .A2 (load_value[9]));
AND2_X4 i_0_0_8 (.ZN (\t_o_values[8] ), .A1 (n_0_0_52), .A2 (load_value[8]));
AND2_X4 i_0_0_7 (.ZN (\t_o_values[7] ), .A1 (n_0_0_52), .A2 (load_value[7]));
AND2_X4 i_0_0_6 (.ZN (\t_o_values[6] ), .A1 (n_0_0_52), .A2 (load_value[6]));
AND2_X1 i_0_0_5 (.ZN (\t_o_values[5] ), .A1 (n_0_0_52), .A2 (load_value[5]));
AND2_X1 i_0_0_4 (.ZN (\t_o_values[4] ), .A1 (n_0_0_52), .A2 (load_value[4]));
AND2_X1 i_0_0_3 (.ZN (\t_o_values[3] ), .A1 (n_0_0_52), .A2 (load_value[3]));
AND2_X1 i_0_0_2 (.ZN (\t_o_values[2] ), .A1 (n_0_0_52), .A2 (load_value[2]));
AND2_X1 i_0_0_1 (.ZN (\t_o_values[1] ), .A1 (n_0_0_52), .A2 (load_value[1]));
AND2_X1 i_0_0_0 (.ZN (\t_o_values[0] ), .A1 (n_0_0_52), .A2 (load_value[0]));
DFF_X1 \o_values_reg[0][0]  (.Q (\o_values[0] [0] ), .CK (n_0_167), .D (sps__n16));
DFF_X1 \o_values_reg[0][1]  (.Q (\o_values[0] [1] ), .CK (n_0_167), .D (sps__n25));
DFF_X1 \o_values_reg[0][2]  (.Q (\o_values[0] [2] ), .CK (n_0_167), .D (sps__n19));
DFF_X1 \o_values_reg[0][3]  (.Q (\o_values[0] [3] ), .CK (n_0_167), .D (sps__n28));
DFF_X1 \o_values_reg[0][4]  (.Q (\o_values[0] [4] ), .CK (n_0_167), .D (sps__n31));
DFF_X1 \o_values_reg[0][5]  (.Q (\o_values[0] [5] ), .CK (n_0_167), .D (sps__n34));
DFF_X1 \o_values_reg[0][6]  (.Q (\o_values[0] [6] ), .CK (n_0_167), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[0][7]  (.Q (\o_values[0] [7] ), .CK (n_0_167), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[0][8]  (.Q (\o_values[0] [8] ), .CK (n_0_167), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[0][9]  (.Q (\o_values[0] [9] ), .CK (n_0_167), .D (sps__n37));
DFF_X1 \o_values_reg[0][10]  (.Q (\o_values[0] [10] ), .CK (n_0_167), .D (sps__n4));
DFF_X1 \o_values_reg[0][11]  (.Q (\o_values[0] [11] ), .CK (n_0_167), .D (sps__n10));
DFF_X1 \o_values_reg[0][12]  (.Q (\o_values[0] [12] ), .CK (n_0_167), .D (sps__n7));
DFF_X1 \o_values_reg[0][13]  (.Q (\o_values[0] [13] ), .CK (n_0_167), .D (sps__n1));
DFF_X1 \o_values_reg[0][14]  (.Q (\o_values[0] [14] ), .CK (n_0_167), .D (sps__n13));
DFF_X1 \o_values_reg[0][15]  (.Q (\o_values[0] [15] ), .CK (n_0_167), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[0]_reg  (.GCK (n_0_167), .CK (clk), .E (n_0_83), .SE (1'b0 ));
DFF_X1 \o_values_reg[1][0]  (.Q (\o_values[1] [0] ), .CK (n_0_166), .D (sps__n16));
DFF_X1 \o_values_reg[1][1]  (.Q (\o_values[1] [1] ), .CK (n_0_166), .D (sps__n25));
DFF_X1 \o_values_reg[1][2]  (.Q (\o_values[1] [2] ), .CK (n_0_166), .D (sps__n19));
DFF_X1 \o_values_reg[1][3]  (.Q (\o_values[1] [3] ), .CK (n_0_166), .D (sps__n28));
DFF_X1 \o_values_reg[1][4]  (.Q (\o_values[1] [4] ), .CK (n_0_166), .D (sps__n31));
DFF_X1 \o_values_reg[1][5]  (.Q (\o_values[1] [5] ), .CK (n_0_166), .D (sps__n34));
DFF_X1 \o_values_reg[1][6]  (.Q (\o_values[1] [6] ), .CK (n_0_166), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[1][7]  (.Q (\o_values[1] [7] ), .CK (n_0_166), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[1][8]  (.Q (\o_values[1] [8] ), .CK (n_0_166), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[1][9]  (.Q (\o_values[1] [9] ), .CK (n_0_166), .D (sps__n37));
DFF_X1 \o_values_reg[1][10]  (.Q (\o_values[1] [10] ), .CK (n_0_166), .D (sps__n4));
DFF_X1 \o_values_reg[1][11]  (.Q (\o_values[1] [11] ), .CK (n_0_166), .D (sps__n10));
DFF_X1 \o_values_reg[1][12]  (.Q (\o_values[1] [12] ), .CK (n_0_166), .D (sps__n7));
DFF_X1 \o_values_reg[1][13]  (.Q (\o_values[1] [13] ), .CK (n_0_166), .D (sps__n1));
DFF_X1 \o_values_reg[1][14]  (.Q (\o_values[1] [14] ), .CK (n_0_166), .D (sps__n13));
DFF_X1 \o_values_reg[1][15]  (.Q (\o_values[1] [15] ), .CK (n_0_166), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[1]_reg  (.GCK (n_0_166), .CK (clk), .E (n_0_82), .SE (1'b0 ));
DFF_X1 \o_values_reg[2][0]  (.Q (\o_values[2] [0] ), .CK (n_0_165), .D (sps__n16));
DFF_X1 \o_values_reg[2][1]  (.Q (\o_values[2] [1] ), .CK (n_0_165), .D (sps__n25));
DFF_X1 \o_values_reg[2][2]  (.Q (\o_values[2] [2] ), .CK (n_0_165), .D (sps__n19));
DFF_X1 \o_values_reg[2][3]  (.Q (\o_values[2] [3] ), .CK (n_0_165), .D (sps__n28));
DFF_X1 \o_values_reg[2][4]  (.Q (\o_values[2] [4] ), .CK (n_0_165), .D (sps__n31));
DFF_X1 \o_values_reg[2][5]  (.Q (\o_values[2] [5] ), .CK (n_0_165), .D (sps__n34));
DFF_X1 \o_values_reg[2][6]  (.Q (\o_values[2] [6] ), .CK (n_0_165), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[2][7]  (.Q (\o_values[2] [7] ), .CK (n_0_165), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[2][8]  (.Q (\o_values[2] [8] ), .CK (n_0_165), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[2][9]  (.Q (\o_values[2] [9] ), .CK (n_0_165), .D (sps__n37));
DFF_X1 \o_values_reg[2][10]  (.Q (\o_values[2] [10] ), .CK (n_0_165), .D (sps__n4));
DFF_X1 \o_values_reg[2][11]  (.Q (\o_values[2] [11] ), .CK (n_0_165), .D (sps__n10));
DFF_X1 \o_values_reg[2][12]  (.Q (\o_values[2] [12] ), .CK (n_0_165), .D (sps__n7));
DFF_X1 \o_values_reg[2][13]  (.Q (\o_values[2] [13] ), .CK (n_0_165), .D (sps__n1));
DFF_X1 \o_values_reg[2][14]  (.Q (\o_values[2] [14] ), .CK (n_0_165), .D (sps__n13));
DFF_X1 \o_values_reg[2][15]  (.Q (\o_values[2] [15] ), .CK (n_0_165), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[2]_reg  (.GCK (n_0_165), .CK (clk), .E (n_0_81), .SE (1'b0 ));
DFF_X1 \o_values_reg[3][0]  (.Q (\o_values[3] [0] ), .CK (n_0_164), .D (sps__n16));
DFF_X1 \o_values_reg[3][1]  (.Q (\o_values[3] [1] ), .CK (n_0_164), .D (sps__n25));
DFF_X1 \o_values_reg[3][2]  (.Q (\o_values[3] [2] ), .CK (n_0_164), .D (sps__n19));
DFF_X1 \o_values_reg[3][3]  (.Q (\o_values[3] [3] ), .CK (n_0_164), .D (sps__n28));
DFF_X1 \o_values_reg[3][4]  (.Q (\o_values[3] [4] ), .CK (n_0_164), .D (sps__n31));
DFF_X1 \o_values_reg[3][5]  (.Q (\o_values[3] [5] ), .CK (n_0_164), .D (sps__n34));
DFF_X1 \o_values_reg[3][6]  (.Q (\o_values[3] [6] ), .CK (n_0_164), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[3][7]  (.Q (\o_values[3] [7] ), .CK (n_0_164), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[3][8]  (.Q (\o_values[3] [8] ), .CK (n_0_164), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[3][9]  (.Q (\o_values[3] [9] ), .CK (n_0_164), .D (sps__n37));
DFF_X1 \o_values_reg[3][10]  (.Q (\o_values[3] [10] ), .CK (n_0_164), .D (sps__n4));
DFF_X1 \o_values_reg[3][11]  (.Q (\o_values[3] [11] ), .CK (n_0_164), .D (sps__n10));
DFF_X1 \o_values_reg[3][12]  (.Q (\o_values[3] [12] ), .CK (n_0_164), .D (sps__n7));
DFF_X1 \o_values_reg[3][13]  (.Q (\o_values[3] [13] ), .CK (n_0_164), .D (sps__n1));
DFF_X1 \o_values_reg[3][14]  (.Q (\o_values[3] [14] ), .CK (n_0_164), .D (sps__n13));
DFF_X1 \o_values_reg[3][15]  (.Q (\o_values[3] [15] ), .CK (n_0_164), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[3]_reg  (.GCK (n_0_164), .CK (clk), .E (n_0_80), .SE (1'b0 ));
DFF_X1 \o_values_reg[4][0]  (.Q (\o_values[4] [0] ), .CK (n_0_163), .D (sps__n16));
DFF_X1 \o_values_reg[4][1]  (.Q (\o_values[4] [1] ), .CK (n_0_163), .D (sps__n25));
DFF_X1 \o_values_reg[4][2]  (.Q (\o_values[4] [2] ), .CK (n_0_163), .D (sps__n19));
DFF_X1 \o_values_reg[4][3]  (.Q (\o_values[4] [3] ), .CK (n_0_163), .D (sps__n28));
DFF_X1 \o_values_reg[4][4]  (.Q (\o_values[4] [4] ), .CK (n_0_163), .D (sps__n31));
DFF_X1 \o_values_reg[4][5]  (.Q (\o_values[4] [5] ), .CK (n_0_163), .D (sps__n34));
DFF_X1 \o_values_reg[4][6]  (.Q (\o_values[4] [6] ), .CK (n_0_163), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[4][7]  (.Q (\o_values[4] [7] ), .CK (n_0_163), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[4][8]  (.Q (\o_values[4] [8] ), .CK (n_0_163), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[4][9]  (.Q (\o_values[4] [9] ), .CK (n_0_163), .D (sps__n37));
DFF_X1 \o_values_reg[4][10]  (.Q (\o_values[4] [10] ), .CK (n_0_163), .D (sps__n4));
DFF_X1 \o_values_reg[4][11]  (.Q (\o_values[4] [11] ), .CK (n_0_163), .D (sps__n10));
DFF_X1 \o_values_reg[4][12]  (.Q (\o_values[4] [12] ), .CK (n_0_163), .D (sps__n7));
DFF_X1 \o_values_reg[4][13]  (.Q (\o_values[4] [13] ), .CK (n_0_163), .D (sps__n1));
DFF_X1 \o_values_reg[4][14]  (.Q (\o_values[4] [14] ), .CK (n_0_163), .D (sps__n13));
DFF_X1 \o_values_reg[4][15]  (.Q (\o_values[4] [15] ), .CK (n_0_163), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[4]_reg  (.GCK (n_0_163), .CK (clk), .E (n_0_79), .SE (1'b0 ));
DFF_X1 \o_values_reg[5][0]  (.Q (\o_values[5] [0] ), .CK (n_0_162), .D (sps__n16));
DFF_X1 \o_values_reg[5][1]  (.Q (\o_values[5] [1] ), .CK (n_0_162), .D (sps__n25));
DFF_X1 \o_values_reg[5][2]  (.Q (\o_values[5] [2] ), .CK (n_0_162), .D (sps__n19));
DFF_X1 \o_values_reg[5][3]  (.Q (\o_values[5] [3] ), .CK (n_0_162), .D (sps__n28));
DFF_X1 \o_values_reg[5][4]  (.Q (\o_values[5] [4] ), .CK (n_0_162), .D (sps__n31));
DFF_X1 \o_values_reg[5][5]  (.Q (\o_values[5] [5] ), .CK (n_0_162), .D (sps__n34));
DFF_X1 \o_values_reg[5][6]  (.Q (\o_values[5] [6] ), .CK (n_0_162), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[5][7]  (.Q (\o_values[5] [7] ), .CK (n_0_162), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[5][8]  (.Q (\o_values[5] [8] ), .CK (n_0_162), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[5][9]  (.Q (\o_values[5] [9] ), .CK (n_0_162), .D (sps__n37));
DFF_X1 \o_values_reg[5][10]  (.Q (\o_values[5] [10] ), .CK (n_0_162), .D (sps__n4));
DFF_X1 \o_values_reg[5][11]  (.Q (\o_values[5] [11] ), .CK (n_0_162), .D (sps__n10));
DFF_X1 \o_values_reg[5][12]  (.Q (\o_values[5] [12] ), .CK (n_0_162), .D (sps__n7));
DFF_X1 \o_values_reg[5][13]  (.Q (\o_values[5] [13] ), .CK (n_0_162), .D (sps__n1));
DFF_X1 \o_values_reg[5][14]  (.Q (\o_values[5] [14] ), .CK (n_0_162), .D (sps__n13));
DFF_X1 \o_values_reg[5][15]  (.Q (\o_values[5] [15] ), .CK (n_0_162), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[5]_reg  (.GCK (n_0_162), .CK (clk), .E (n_0_78), .SE (1'b0 ));
DFF_X1 \o_values_reg[6][0]  (.Q (\o_values[6] [0] ), .CK (n_0_161), .D (sps__n16));
DFF_X1 \o_values_reg[6][1]  (.Q (\o_values[6] [1] ), .CK (n_0_161), .D (sps__n25));
DFF_X1 \o_values_reg[6][2]  (.Q (\o_values[6] [2] ), .CK (n_0_161), .D (sps__n19));
DFF_X1 \o_values_reg[6][3]  (.Q (\o_values[6] [3] ), .CK (n_0_161), .D (sps__n28));
DFF_X1 \o_values_reg[6][4]  (.Q (\o_values[6] [4] ), .CK (n_0_161), .D (sps__n31));
DFF_X1 \o_values_reg[6][5]  (.Q (\o_values[6] [5] ), .CK (n_0_161), .D (sps__n34));
DFF_X1 \o_values_reg[6][6]  (.Q (\o_values[6] [6] ), .CK (n_0_161), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[6][7]  (.Q (\o_values[6] [7] ), .CK (n_0_161), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[6][8]  (.Q (\o_values[6] [8] ), .CK (n_0_161), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[6][9]  (.Q (\o_values[6] [9] ), .CK (n_0_161), .D (sps__n37));
DFF_X1 \o_values_reg[6][10]  (.Q (\o_values[6] [10] ), .CK (n_0_161), .D (sps__n4));
DFF_X1 \o_values_reg[6][11]  (.Q (\o_values[6] [11] ), .CK (n_0_161), .D (sps__n10));
DFF_X1 \o_values_reg[6][12]  (.Q (\o_values[6] [12] ), .CK (n_0_161), .D (sps__n7));
DFF_X1 \o_values_reg[6][13]  (.Q (\o_values[6] [13] ), .CK (n_0_161), .D (sps__n1));
DFF_X1 \o_values_reg[6][14]  (.Q (\o_values[6] [14] ), .CK (n_0_161), .D (sps__n13));
DFF_X1 \o_values_reg[6][15]  (.Q (\o_values[6] [15] ), .CK (n_0_161), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[6]_reg  (.GCK (n_0_161), .CK (clk), .E (n_0_77), .SE (1'b0 ));
DFF_X1 \o_values_reg[7][0]  (.Q (\o_values[7] [0] ), .CK (n_0_160), .D (sps__n16));
DFF_X1 \o_values_reg[7][1]  (.Q (\o_values[7] [1] ), .CK (n_0_160), .D (sps__n25));
DFF_X1 \o_values_reg[7][2]  (.Q (\o_values[7] [2] ), .CK (n_0_160), .D (sps__n19));
DFF_X1 \o_values_reg[7][3]  (.Q (\o_values[7] [3] ), .CK (n_0_160), .D (sps__n28));
DFF_X1 \o_values_reg[7][4]  (.Q (\o_values[7] [4] ), .CK (n_0_160), .D (sps__n31));
DFF_X1 \o_values_reg[7][5]  (.Q (\o_values[7] [5] ), .CK (n_0_160), .D (sps__n34));
DFF_X1 \o_values_reg[7][6]  (.Q (\o_values[7] [6] ), .CK (n_0_160), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[7][7]  (.Q (\o_values[7] [7] ), .CK (n_0_160), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[7][8]  (.Q (\o_values[7] [8] ), .CK (n_0_160), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[7][9]  (.Q (\o_values[7] [9] ), .CK (n_0_160), .D (sps__n37));
DFF_X1 \o_values_reg[7][10]  (.Q (\o_values[7] [10] ), .CK (n_0_160), .D (sps__n4));
DFF_X1 \o_values_reg[7][11]  (.Q (\o_values[7] [11] ), .CK (n_0_160), .D (sps__n10));
DFF_X1 \o_values_reg[7][12]  (.Q (\o_values[7] [12] ), .CK (n_0_160), .D (sps__n7));
DFF_X1 \o_values_reg[7][13]  (.Q (\o_values[7] [13] ), .CK (n_0_160), .D (sps__n1));
DFF_X1 \o_values_reg[7][14]  (.Q (\o_values[7] [14] ), .CK (n_0_160), .D (sps__n13));
DFF_X1 \o_values_reg[7][15]  (.Q (\o_values[7] [15] ), .CK (n_0_160), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[7]_reg  (.GCK (n_0_160), .CK (clk), .E (n_0_76), .SE (1'b0 ));
DFF_X1 \o_values_reg[8][0]  (.Q (\o_values[8] [0] ), .CK (n_0_159), .D (sps__n16));
DFF_X1 \o_values_reg[8][1]  (.Q (\o_values[8] [1] ), .CK (n_0_159), .D (sps__n25));
DFF_X1 \o_values_reg[8][2]  (.Q (\o_values[8] [2] ), .CK (n_0_159), .D (sps__n19));
DFF_X1 \o_values_reg[8][3]  (.Q (\o_values[8] [3] ), .CK (n_0_159), .D (sps__n28));
DFF_X1 \o_values_reg[8][4]  (.Q (\o_values[8] [4] ), .CK (n_0_159), .D (sps__n31));
DFF_X1 \o_values_reg[8][5]  (.Q (\o_values[8] [5] ), .CK (n_0_159), .D (sps__n34));
DFF_X1 \o_values_reg[8][6]  (.Q (\o_values[8] [6] ), .CK (n_0_159), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[8][7]  (.Q (\o_values[8] [7] ), .CK (n_0_159), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[8][8]  (.Q (\o_values[8] [8] ), .CK (n_0_159), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[8][9]  (.Q (\o_values[8] [9] ), .CK (n_0_159), .D (sps__n37));
DFF_X1 \o_values_reg[8][10]  (.Q (\o_values[8] [10] ), .CK (n_0_159), .D (sps__n4));
DFF_X1 \o_values_reg[8][11]  (.Q (\o_values[8] [11] ), .CK (n_0_159), .D (sps__n10));
DFF_X1 \o_values_reg[8][12]  (.Q (\o_values[8] [12] ), .CK (n_0_159), .D (sps__n7));
DFF_X1 \o_values_reg[8][13]  (.Q (\o_values[8] [13] ), .CK (n_0_159), .D (sps__n1));
DFF_X1 \o_values_reg[8][14]  (.Q (\o_values[8] [14] ), .CK (n_0_159), .D (sps__n13));
DFF_X1 \o_values_reg[8][15]  (.Q (\o_values[8] [15] ), .CK (n_0_159), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[8]_reg  (.GCK (n_0_159), .CK (clk), .E (n_0_75), .SE (1'b0 ));
DFF_X1 \o_values_reg[9][0]  (.Q (\o_values[9] [0] ), .CK (n_0_158), .D (sps__n16));
DFF_X1 \o_values_reg[9][1]  (.Q (\o_values[9] [1] ), .CK (n_0_158), .D (sps__n25));
DFF_X1 \o_values_reg[9][2]  (.Q (\o_values[9] [2] ), .CK (n_0_158), .D (sps__n19));
DFF_X1 \o_values_reg[9][3]  (.Q (\o_values[9] [3] ), .CK (n_0_158), .D (sps__n28));
DFF_X1 \o_values_reg[9][4]  (.Q (\o_values[9] [4] ), .CK (n_0_158), .D (sps__n31));
DFF_X1 \o_values_reg[9][5]  (.Q (\o_values[9] [5] ), .CK (n_0_158), .D (sps__n34));
DFF_X1 \o_values_reg[9][6]  (.Q (\o_values[9] [6] ), .CK (n_0_158), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[9][7]  (.Q (\o_values[9] [7] ), .CK (n_0_158), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[9][8]  (.Q (\o_values[9] [8] ), .CK (n_0_158), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[9][9]  (.Q (\o_values[9] [9] ), .CK (n_0_158), .D (sps__n37));
DFF_X1 \o_values_reg[9][10]  (.Q (\o_values[9] [10] ), .CK (n_0_158), .D (sps__n4));
DFF_X1 \o_values_reg[9][11]  (.Q (\o_values[9] [11] ), .CK (n_0_158), .D (sps__n10));
DFF_X1 \o_values_reg[9][12]  (.Q (\o_values[9] [12] ), .CK (n_0_158), .D (sps__n7));
DFF_X1 \o_values_reg[9][13]  (.Q (\o_values[9] [13] ), .CK (n_0_158), .D (sps__n1));
DFF_X1 \o_values_reg[9][14]  (.Q (\o_values[9] [14] ), .CK (n_0_158), .D (sps__n13));
DFF_X1 \o_values_reg[9][15]  (.Q (\o_values[9] [15] ), .CK (n_0_158), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[9]_reg  (.GCK (n_0_158), .CK (clk), .E (n_0_74), .SE (1'b0 ));
DFF_X1 \o_values_reg[10][0]  (.Q (\o_values[10] [0] ), .CK (n_0_157), .D (sps__n16));
DFF_X1 \o_values_reg[10][1]  (.Q (\o_values[10] [1] ), .CK (n_0_157), .D (sps__n25));
DFF_X1 \o_values_reg[10][2]  (.Q (\o_values[10] [2] ), .CK (n_0_157), .D (sps__n19));
DFF_X1 \o_values_reg[10][3]  (.Q (\o_values[10] [3] ), .CK (n_0_157), .D (sps__n28));
DFF_X1 \o_values_reg[10][4]  (.Q (\o_values[10] [4] ), .CK (n_0_157), .D (sps__n31));
DFF_X1 \o_values_reg[10][5]  (.Q (\o_values[10] [5] ), .CK (n_0_157), .D (sps__n34));
DFF_X1 \o_values_reg[10][6]  (.Q (\o_values[10] [6] ), .CK (n_0_157), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[10][7]  (.Q (\o_values[10] [7] ), .CK (n_0_157), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[10][8]  (.Q (\o_values[10] [8] ), .CK (n_0_157), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[10][9]  (.Q (\o_values[10] [9] ), .CK (n_0_157), .D (sps__n37));
DFF_X1 \o_values_reg[10][10]  (.Q (\o_values[10] [10] ), .CK (n_0_157), .D (sps__n4));
DFF_X1 \o_values_reg[10][11]  (.Q (\o_values[10] [11] ), .CK (n_0_157), .D (sps__n10));
DFF_X1 \o_values_reg[10][12]  (.Q (\o_values[10] [12] ), .CK (n_0_157), .D (sps__n7));
DFF_X1 \o_values_reg[10][13]  (.Q (\o_values[10] [13] ), .CK (n_0_157), .D (sps__n1));
DFF_X1 \o_values_reg[10][14]  (.Q (\o_values[10] [14] ), .CK (n_0_157), .D (sps__n13));
DFF_X1 \o_values_reg[10][15]  (.Q (\o_values[10] [15] ), .CK (n_0_157), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[10]_reg  (.GCK (n_0_157), .CK (clk), .E (n_0_73), .SE (1'b0 ));
DFF_X1 \o_values_reg[11][0]  (.Q (\o_values[11] [0] ), .CK (n_0_156), .D (sps__n16));
DFF_X1 \o_values_reg[11][1]  (.Q (\o_values[11] [1] ), .CK (n_0_156), .D (sps__n25));
DFF_X1 \o_values_reg[11][2]  (.Q (\o_values[11] [2] ), .CK (n_0_156), .D (sps__n19));
DFF_X1 \o_values_reg[11][3]  (.Q (\o_values[11] [3] ), .CK (n_0_156), .D (sps__n28));
DFF_X1 \o_values_reg[11][4]  (.Q (\o_values[11] [4] ), .CK (n_0_156), .D (sps__n31));
DFF_X1 \o_values_reg[11][5]  (.Q (\o_values[11] [5] ), .CK (n_0_156), .D (sps__n34));
DFF_X1 \o_values_reg[11][6]  (.Q (\o_values[11] [6] ), .CK (n_0_156), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[11][7]  (.Q (\o_values[11] [7] ), .CK (n_0_156), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[11][8]  (.Q (\o_values[11] [8] ), .CK (n_0_156), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[11][9]  (.Q (\o_values[11] [9] ), .CK (n_0_156), .D (sps__n37));
DFF_X1 \o_values_reg[11][10]  (.Q (\o_values[11] [10] ), .CK (n_0_156), .D (sps__n4));
DFF_X1 \o_values_reg[11][11]  (.Q (\o_values[11] [11] ), .CK (n_0_156), .D (sps__n10));
DFF_X1 \o_values_reg[11][12]  (.Q (\o_values[11] [12] ), .CK (n_0_156), .D (sps__n7));
DFF_X1 \o_values_reg[11][13]  (.Q (\o_values[11] [13] ), .CK (n_0_156), .D (sps__n1));
DFF_X1 \o_values_reg[11][14]  (.Q (\o_values[11] [14] ), .CK (n_0_156), .D (sps__n13));
DFF_X1 \o_values_reg[11][15]  (.Q (\o_values[11] [15] ), .CK (n_0_156), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[11]_reg  (.GCK (n_0_156), .CK (clk), .E (n_0_72), .SE (1'b0 ));
DFF_X1 \o_values_reg[12][0]  (.Q (\o_values[12] [0] ), .CK (n_0_155), .D (sps__n16));
DFF_X1 \o_values_reg[12][1]  (.Q (\o_values[12] [1] ), .CK (n_0_155), .D (sps__n25));
DFF_X1 \o_values_reg[12][2]  (.Q (\o_values[12] [2] ), .CK (n_0_155), .D (sps__n19));
DFF_X1 \o_values_reg[12][3]  (.Q (\o_values[12] [3] ), .CK (n_0_155), .D (sps__n28));
DFF_X1 \o_values_reg[12][4]  (.Q (\o_values[12] [4] ), .CK (n_0_155), .D (sps__n31));
DFF_X1 \o_values_reg[12][5]  (.Q (\o_values[12] [5] ), .CK (n_0_155), .D (sps__n34));
DFF_X1 \o_values_reg[12][6]  (.Q (\o_values[12] [6] ), .CK (n_0_155), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[12][7]  (.Q (\o_values[12] [7] ), .CK (n_0_155), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[12][8]  (.Q (\o_values[12] [8] ), .CK (n_0_155), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[12][9]  (.Q (\o_values[12] [9] ), .CK (n_0_155), .D (sps__n37));
DFF_X1 \o_values_reg[12][10]  (.Q (\o_values[12] [10] ), .CK (n_0_155), .D (sps__n4));
DFF_X1 \o_values_reg[12][11]  (.Q (\o_values[12] [11] ), .CK (n_0_155), .D (sps__n10));
DFF_X1 \o_values_reg[12][12]  (.Q (\o_values[12] [12] ), .CK (n_0_155), .D (sps__n7));
DFF_X1 \o_values_reg[12][13]  (.Q (\o_values[12] [13] ), .CK (n_0_155), .D (sps__n1));
DFF_X1 \o_values_reg[12][14]  (.Q (\o_values[12] [14] ), .CK (n_0_155), .D (sps__n13));
DFF_X1 \o_values_reg[12][15]  (.Q (\o_values[12] [15] ), .CK (n_0_155), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[12]_reg  (.GCK (n_0_155), .CK (clk), .E (n_0_71), .SE (1'b0 ));
DFF_X1 \o_values_reg[13][0]  (.Q (\o_values[13] [0] ), .CK (n_0_154), .D (sps__n16));
DFF_X1 \o_values_reg[13][1]  (.Q (\o_values[13] [1] ), .CK (n_0_154), .D (sps__n25));
DFF_X1 \o_values_reg[13][2]  (.Q (\o_values[13] [2] ), .CK (n_0_154), .D (sps__n19));
DFF_X1 \o_values_reg[13][3]  (.Q (\o_values[13] [3] ), .CK (n_0_154), .D (sps__n28));
DFF_X1 \o_values_reg[13][4]  (.Q (\o_values[13] [4] ), .CK (n_0_154), .D (sps__n31));
DFF_X1 \o_values_reg[13][5]  (.Q (\o_values[13] [5] ), .CK (n_0_154), .D (sps__n34));
DFF_X1 \o_values_reg[13][6]  (.Q (\o_values[13] [6] ), .CK (n_0_154), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[13][7]  (.Q (\o_values[13] [7] ), .CK (n_0_154), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[13][8]  (.Q (\o_values[13] [8] ), .CK (n_0_154), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[13][9]  (.Q (\o_values[13] [9] ), .CK (n_0_154), .D (sps__n37));
DFF_X1 \o_values_reg[13][10]  (.Q (\o_values[13] [10] ), .CK (n_0_154), .D (sps__n4));
DFF_X1 \o_values_reg[13][11]  (.Q (\o_values[13] [11] ), .CK (n_0_154), .D (sps__n10));
DFF_X1 \o_values_reg[13][12]  (.Q (\o_values[13] [12] ), .CK (n_0_154), .D (sps__n7));
DFF_X1 \o_values_reg[13][13]  (.Q (\o_values[13] [13] ), .CK (n_0_154), .D (sps__n1));
DFF_X1 \o_values_reg[13][14]  (.Q (\o_values[13] [14] ), .CK (n_0_154), .D (sps__n13));
DFF_X1 \o_values_reg[13][15]  (.Q (\o_values[13] [15] ), .CK (n_0_154), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[13]_reg  (.GCK (n_0_154), .CK (clk), .E (n_0_70), .SE (1'b0 ));
DFF_X1 \o_values_reg[14][0]  (.Q (\o_values[14] [0] ), .CK (n_0_153), .D (sps__n16));
DFF_X1 \o_values_reg[14][1]  (.Q (\o_values[14] [1] ), .CK (n_0_153), .D (sps__n25));
DFF_X1 \o_values_reg[14][2]  (.Q (\o_values[14] [2] ), .CK (n_0_153), .D (sps__n19));
DFF_X1 \o_values_reg[14][3]  (.Q (\o_values[14] [3] ), .CK (n_0_153), .D (sps__n28));
DFF_X1 \o_values_reg[14][4]  (.Q (\o_values[14] [4] ), .CK (n_0_153), .D (sps__n31));
DFF_X1 \o_values_reg[14][5]  (.Q (\o_values[14] [5] ), .CK (n_0_153), .D (sps__n34));
DFF_X1 \o_values_reg[14][6]  (.Q (\o_values[14] [6] ), .CK (n_0_153), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[14][7]  (.Q (\o_values[14] [7] ), .CK (n_0_153), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[14][8]  (.Q (\o_values[14] [8] ), .CK (n_0_153), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[14][9]  (.Q (\o_values[14] [9] ), .CK (n_0_153), .D (sps__n37));
DFF_X1 \o_values_reg[14][10]  (.Q (\o_values[14] [10] ), .CK (n_0_153), .D (sps__n4));
DFF_X1 \o_values_reg[14][11]  (.Q (\o_values[14] [11] ), .CK (n_0_153), .D (sps__n10));
DFF_X1 \o_values_reg[14][12]  (.Q (\o_values[14] [12] ), .CK (n_0_153), .D (sps__n7));
DFF_X1 \o_values_reg[14][13]  (.Q (\o_values[14] [13] ), .CK (n_0_153), .D (sps__n1));
DFF_X1 \o_values_reg[14][14]  (.Q (\o_values[14] [14] ), .CK (n_0_153), .D (sps__n13));
DFF_X1 \o_values_reg[14][15]  (.Q (\o_values[14] [15] ), .CK (n_0_153), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[14]_reg  (.GCK (n_0_153), .CK (clk), .E (n_0_69), .SE (1'b0 ));
DFF_X1 \o_values_reg[15][0]  (.Q (\o_values[15] [0] ), .CK (n_0_152), .D (sps__n16));
DFF_X1 \o_values_reg[15][1]  (.Q (\o_values[15] [1] ), .CK (n_0_152), .D (sps__n25));
DFF_X1 \o_values_reg[15][2]  (.Q (\o_values[15] [2] ), .CK (n_0_152), .D (sps__n19));
DFF_X1 \o_values_reg[15][3]  (.Q (\o_values[15] [3] ), .CK (n_0_152), .D (sps__n28));
DFF_X1 \o_values_reg[15][4]  (.Q (\o_values[15] [4] ), .CK (n_0_152), .D (sps__n31));
DFF_X1 \o_values_reg[15][5]  (.Q (\o_values[15] [5] ), .CK (n_0_152), .D (sps__n34));
DFF_X1 \o_values_reg[15][6]  (.Q (\o_values[15] [6] ), .CK (n_0_152), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[15][7]  (.Q (\o_values[15] [7] ), .CK (n_0_152), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[15][8]  (.Q (\o_values[15] [8] ), .CK (n_0_152), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[15][9]  (.Q (\o_values[15] [9] ), .CK (n_0_152), .D (sps__n37));
DFF_X1 \o_values_reg[15][10]  (.Q (\o_values[15] [10] ), .CK (n_0_152), .D (sps__n4));
DFF_X1 \o_values_reg[15][11]  (.Q (\o_values[15] [11] ), .CK (n_0_152), .D (sps__n10));
DFF_X1 \o_values_reg[15][12]  (.Q (\o_values[15] [12] ), .CK (n_0_152), .D (sps__n7));
DFF_X1 \o_values_reg[15][13]  (.Q (\o_values[15] [13] ), .CK (n_0_152), .D (sps__n1));
DFF_X1 \o_values_reg[15][14]  (.Q (\o_values[15] [14] ), .CK (n_0_152), .D (sps__n13));
DFF_X1 \o_values_reg[15][15]  (.Q (\o_values[15] [15] ), .CK (n_0_152), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[15]_reg  (.GCK (n_0_152), .CK (clk), .E (n_0_68), .SE (1'b0 ));
DFF_X1 \o_values_reg[16][0]  (.Q (\o_values[16] [0] ), .CK (n_0_151), .D (sps__n16));
DFF_X1 \o_values_reg[16][1]  (.Q (\o_values[16] [1] ), .CK (n_0_151), .D (sps__n25));
DFF_X1 \o_values_reg[16][2]  (.Q (\o_values[16] [2] ), .CK (n_0_151), .D (sps__n19));
DFF_X1 \o_values_reg[16][3]  (.Q (\o_values[16] [3] ), .CK (n_0_151), .D (sps__n28));
DFF_X1 \o_values_reg[16][4]  (.Q (\o_values[16] [4] ), .CK (n_0_151), .D (sps__n31));
DFF_X1 \o_values_reg[16][5]  (.Q (\o_values[16] [5] ), .CK (n_0_151), .D (sps__n34));
DFF_X1 \o_values_reg[16][6]  (.Q (\o_values[16] [6] ), .CK (n_0_151), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[16][7]  (.Q (\o_values[16] [7] ), .CK (n_0_151), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[16][8]  (.Q (\o_values[16] [8] ), .CK (n_0_151), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[16][9]  (.Q (\o_values[16] [9] ), .CK (n_0_151), .D (sps__n37));
DFF_X1 \o_values_reg[16][10]  (.Q (\o_values[16] [10] ), .CK (n_0_151), .D (sps__n4));
DFF_X1 \o_values_reg[16][11]  (.Q (\o_values[16] [11] ), .CK (n_0_151), .D (sps__n10));
DFF_X1 \o_values_reg[16][12]  (.Q (\o_values[16] [12] ), .CK (n_0_151), .D (sps__n7));
DFF_X1 \o_values_reg[16][13]  (.Q (\o_values[16] [13] ), .CK (n_0_151), .D (sps__n1));
DFF_X1 \o_values_reg[16][14]  (.Q (\o_values[16] [14] ), .CK (n_0_151), .D (sps__n13));
DFF_X1 \o_values_reg[16][15]  (.Q (\o_values[16] [15] ), .CK (n_0_151), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[16]_reg  (.GCK (n_0_151), .CK (clk), .E (n_0_67), .SE (1'b0 ));
DFF_X1 \o_values_reg[17][0]  (.Q (\o_values[17] [0] ), .CK (n_0_150), .D (sps__n16));
DFF_X1 \o_values_reg[17][1]  (.Q (\o_values[17] [1] ), .CK (n_0_150), .D (sps__n25));
DFF_X1 \o_values_reg[17][2]  (.Q (\o_values[17] [2] ), .CK (n_0_150), .D (sps__n19));
DFF_X1 \o_values_reg[17][3]  (.Q (\o_values[17] [3] ), .CK (n_0_150), .D (sps__n28));
DFF_X1 \o_values_reg[17][4]  (.Q (\o_values[17] [4] ), .CK (n_0_150), .D (sps__n31));
DFF_X1 \o_values_reg[17][5]  (.Q (\o_values[17] [5] ), .CK (n_0_150), .D (sps__n34));
DFF_X1 \o_values_reg[17][6]  (.Q (\o_values[17] [6] ), .CK (n_0_150), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[17][7]  (.Q (\o_values[17] [7] ), .CK (n_0_150), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[17][8]  (.Q (\o_values[17] [8] ), .CK (n_0_150), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[17][9]  (.Q (\o_values[17] [9] ), .CK (n_0_150), .D (sps__n37));
DFF_X1 \o_values_reg[17][10]  (.Q (\o_values[17] [10] ), .CK (n_0_150), .D (sps__n4));
DFF_X1 \o_values_reg[17][11]  (.Q (\o_values[17] [11] ), .CK (n_0_150), .D (sps__n10));
DFF_X1 \o_values_reg[17][12]  (.Q (\o_values[17] [12] ), .CK (n_0_150), .D (sps__n7));
DFF_X1 \o_values_reg[17][13]  (.Q (\o_values[17] [13] ), .CK (n_0_150), .D (sps__n1));
DFF_X1 \o_values_reg[17][14]  (.Q (\o_values[17] [14] ), .CK (n_0_150), .D (sps__n13));
DFF_X1 \o_values_reg[17][15]  (.Q (\o_values[17] [15] ), .CK (n_0_150), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[17]_reg  (.GCK (n_0_150), .CK (clk), .E (n_0_66), .SE (1'b0 ));
DFF_X1 \o_values_reg[18][0]  (.Q (\o_values[18] [0] ), .CK (n_0_149), .D (sps__n16));
DFF_X1 \o_values_reg[18][1]  (.Q (\o_values[18] [1] ), .CK (n_0_149), .D (sps__n25));
DFF_X1 \o_values_reg[18][2]  (.Q (\o_values[18] [2] ), .CK (n_0_149), .D (sps__n19));
DFF_X1 \o_values_reg[18][3]  (.Q (\o_values[18] [3] ), .CK (n_0_149), .D (sps__n28));
DFF_X1 \o_values_reg[18][4]  (.Q (\o_values[18] [4] ), .CK (n_0_149), .D (sps__n31));
DFF_X1 \o_values_reg[18][5]  (.Q (\o_values[18] [5] ), .CK (n_0_149), .D (sps__n34));
DFF_X1 \o_values_reg[18][6]  (.Q (\o_values[18] [6] ), .CK (n_0_149), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[18][7]  (.Q (\o_values[18] [7] ), .CK (n_0_149), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[18][8]  (.Q (\o_values[18] [8] ), .CK (n_0_149), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[18][9]  (.Q (\o_values[18] [9] ), .CK (n_0_149), .D (sps__n37));
DFF_X1 \o_values_reg[18][10]  (.Q (\o_values[18] [10] ), .CK (n_0_149), .D (sps__n4));
DFF_X1 \o_values_reg[18][11]  (.Q (\o_values[18] [11] ), .CK (n_0_149), .D (sps__n10));
DFF_X1 \o_values_reg[18][12]  (.Q (\o_values[18] [12] ), .CK (n_0_149), .D (sps__n7));
DFF_X1 \o_values_reg[18][13]  (.Q (\o_values[18] [13] ), .CK (n_0_149), .D (sps__n1));
DFF_X1 \o_values_reg[18][14]  (.Q (\o_values[18] [14] ), .CK (n_0_149), .D (sps__n13));
DFF_X1 \o_values_reg[18][15]  (.Q (\o_values[18] [15] ), .CK (n_0_149), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[18]_reg  (.GCK (n_0_149), .CK (clk), .E (n_0_65), .SE (1'b0 ));
DFF_X1 \o_values_reg[19][0]  (.Q (\o_values[19] [0] ), .CK (n_0_148), .D (sps__n16));
DFF_X1 \o_values_reg[19][1]  (.Q (\o_values[19] [1] ), .CK (n_0_148), .D (sps__n25));
DFF_X1 \o_values_reg[19][2]  (.Q (\o_values[19] [2] ), .CK (n_0_148), .D (sps__n19));
DFF_X1 \o_values_reg[19][3]  (.Q (\o_values[19] [3] ), .CK (n_0_148), .D (sps__n28));
DFF_X1 \o_values_reg[19][4]  (.Q (\o_values[19] [4] ), .CK (n_0_148), .D (sps__n31));
DFF_X1 \o_values_reg[19][5]  (.Q (\o_values[19] [5] ), .CK (n_0_148), .D (sps__n34));
DFF_X1 \o_values_reg[19][6]  (.Q (\o_values[19] [6] ), .CK (n_0_148), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[19][7]  (.Q (\o_values[19] [7] ), .CK (n_0_148), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[19][8]  (.Q (\o_values[19] [8] ), .CK (n_0_148), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[19][9]  (.Q (\o_values[19] [9] ), .CK (n_0_148), .D (sps__n37));
DFF_X1 \o_values_reg[19][10]  (.Q (\o_values[19] [10] ), .CK (n_0_148), .D (sps__n4));
DFF_X1 \o_values_reg[19][11]  (.Q (\o_values[19] [11] ), .CK (n_0_148), .D (sps__n10));
DFF_X1 \o_values_reg[19][12]  (.Q (\o_values[19] [12] ), .CK (n_0_148), .D (sps__n7));
DFF_X1 \o_values_reg[19][13]  (.Q (\o_values[19] [13] ), .CK (n_0_148), .D (sps__n1));
DFF_X1 \o_values_reg[19][14]  (.Q (\o_values[19] [14] ), .CK (n_0_148), .D (sps__n13));
DFF_X1 \o_values_reg[19][15]  (.Q (\o_values[19] [15] ), .CK (n_0_148), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[19]_reg  (.GCK (n_0_148), .CK (clk), .E (n_0_64), .SE (1'b0 ));
DFF_X1 \o_values_reg[20][0]  (.Q (\o_values[20] [0] ), .CK (n_0_147), .D (sps__n16));
DFF_X1 \o_values_reg[20][1]  (.Q (\o_values[20] [1] ), .CK (n_0_147), .D (sps__n25));
DFF_X1 \o_values_reg[20][2]  (.Q (\o_values[20] [2] ), .CK (n_0_147), .D (sps__n19));
DFF_X1 \o_values_reg[20][3]  (.Q (\o_values[20] [3] ), .CK (n_0_147), .D (sps__n28));
DFF_X1 \o_values_reg[20][4]  (.Q (\o_values[20] [4] ), .CK (n_0_147), .D (sps__n31));
DFF_X1 \o_values_reg[20][5]  (.Q (\o_values[20] [5] ), .CK (n_0_147), .D (sps__n34));
DFF_X1 \o_values_reg[20][6]  (.Q (\o_values[20] [6] ), .CK (n_0_147), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[20][7]  (.Q (\o_values[20] [7] ), .CK (n_0_147), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[20][8]  (.Q (\o_values[20] [8] ), .CK (n_0_147), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[20][9]  (.Q (\o_values[20] [9] ), .CK (n_0_147), .D (sps__n37));
DFF_X1 \o_values_reg[20][10]  (.Q (\o_values[20] [10] ), .CK (n_0_147), .D (sps__n4));
DFF_X1 \o_values_reg[20][11]  (.Q (\o_values[20] [11] ), .CK (n_0_147), .D (sps__n10));
DFF_X1 \o_values_reg[20][12]  (.Q (\o_values[20] [12] ), .CK (n_0_147), .D (sps__n7));
DFF_X1 \o_values_reg[20][13]  (.Q (\o_values[20] [13] ), .CK (n_0_147), .D (sps__n1));
DFF_X1 \o_values_reg[20][14]  (.Q (\o_values[20] [14] ), .CK (n_0_147), .D (sps__n13));
DFF_X1 \o_values_reg[20][15]  (.Q (\o_values[20] [15] ), .CK (n_0_147), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[20]_reg  (.GCK (n_0_147), .CK (clk), .E (n_0_63), .SE (1'b0 ));
DFF_X1 \o_values_reg[21][0]  (.Q (\o_values[21] [0] ), .CK (n_0_146), .D (sps__n16));
DFF_X1 \o_values_reg[21][1]  (.Q (\o_values[21] [1] ), .CK (n_0_146), .D (sps__n25));
DFF_X1 \o_values_reg[21][2]  (.Q (\o_values[21] [2] ), .CK (n_0_146), .D (sps__n19));
DFF_X1 \o_values_reg[21][3]  (.Q (\o_values[21] [3] ), .CK (n_0_146), .D (sps__n28));
DFF_X1 \o_values_reg[21][4]  (.Q (\o_values[21] [4] ), .CK (n_0_146), .D (sps__n31));
DFF_X1 \o_values_reg[21][5]  (.Q (\o_values[21] [5] ), .CK (n_0_146), .D (sps__n34));
DFF_X1 \o_values_reg[21][6]  (.Q (\o_values[21] [6] ), .CK (n_0_146), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[21][7]  (.Q (\o_values[21] [7] ), .CK (n_0_146), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[21][8]  (.Q (\o_values[21] [8] ), .CK (n_0_146), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[21][9]  (.Q (\o_values[21] [9] ), .CK (n_0_146), .D (sps__n37));
DFF_X1 \o_values_reg[21][10]  (.Q (\o_values[21] [10] ), .CK (n_0_146), .D (sps__n4));
DFF_X1 \o_values_reg[21][11]  (.Q (\o_values[21] [11] ), .CK (n_0_146), .D (sps__n10));
DFF_X1 \o_values_reg[21][12]  (.Q (\o_values[21] [12] ), .CK (n_0_146), .D (sps__n7));
DFF_X1 \o_values_reg[21][13]  (.Q (\o_values[21] [13] ), .CK (n_0_146), .D (sps__n1));
DFF_X1 \o_values_reg[21][14]  (.Q (\o_values[21] [14] ), .CK (n_0_146), .D (sps__n13));
DFF_X1 \o_values_reg[21][15]  (.Q (\o_values[21] [15] ), .CK (n_0_146), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[21]_reg  (.GCK (n_0_146), .CK (clk), .E (n_0_62), .SE (1'b0 ));
DFF_X1 \o_values_reg[22][0]  (.Q (\o_values[22] [0] ), .CK (n_0_145), .D (sps__n16));
DFF_X1 \o_values_reg[22][1]  (.Q (\o_values[22] [1] ), .CK (n_0_145), .D (sps__n25));
DFF_X1 \o_values_reg[22][2]  (.Q (\o_values[22] [2] ), .CK (n_0_145), .D (sps__n19));
DFF_X1 \o_values_reg[22][3]  (.Q (\o_values[22] [3] ), .CK (n_0_145), .D (sps__n28));
DFF_X1 \o_values_reg[22][4]  (.Q (\o_values[22] [4] ), .CK (n_0_145), .D (sps__n31));
DFF_X1 \o_values_reg[22][5]  (.Q (\o_values[22] [5] ), .CK (n_0_145), .D (sps__n34));
DFF_X1 \o_values_reg[22][6]  (.Q (\o_values[22] [6] ), .CK (n_0_145), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[22][7]  (.Q (\o_values[22] [7] ), .CK (n_0_145), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[22][8]  (.Q (\o_values[22] [8] ), .CK (n_0_145), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[22][9]  (.Q (\o_values[22] [9] ), .CK (n_0_145), .D (sps__n37));
DFF_X1 \o_values_reg[22][10]  (.Q (\o_values[22] [10] ), .CK (n_0_145), .D (sps__n4));
DFF_X1 \o_values_reg[22][11]  (.Q (\o_values[22] [11] ), .CK (n_0_145), .D (sps__n10));
DFF_X1 \o_values_reg[22][12]  (.Q (\o_values[22] [12] ), .CK (n_0_145), .D (sps__n7));
DFF_X1 \o_values_reg[22][13]  (.Q (\o_values[22] [13] ), .CK (n_0_145), .D (sps__n1));
DFF_X1 \o_values_reg[22][14]  (.Q (\o_values[22] [14] ), .CK (n_0_145), .D (sps__n13));
DFF_X1 \o_values_reg[22][15]  (.Q (\o_values[22] [15] ), .CK (n_0_145), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[22]_reg  (.GCK (n_0_145), .CK (clk), .E (n_0_61), .SE (1'b0 ));
DFF_X1 \o_values_reg[23][0]  (.Q (\o_values[23] [0] ), .CK (n_0_144), .D (sps__n16));
DFF_X1 \o_values_reg[23][1]  (.Q (\o_values[23] [1] ), .CK (n_0_144), .D (sps__n25));
DFF_X1 \o_values_reg[23][2]  (.Q (\o_values[23] [2] ), .CK (n_0_144), .D (sps__n19));
DFF_X1 \o_values_reg[23][3]  (.Q (\o_values[23] [3] ), .CK (n_0_144), .D (sps__n28));
DFF_X1 \o_values_reg[23][4]  (.Q (\o_values[23] [4] ), .CK (n_0_144), .D (sps__n31));
DFF_X1 \o_values_reg[23][5]  (.Q (\o_values[23] [5] ), .CK (n_0_144), .D (sps__n34));
DFF_X1 \o_values_reg[23][6]  (.Q (\o_values[23] [6] ), .CK (n_0_144), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[23][7]  (.Q (\o_values[23] [7] ), .CK (n_0_144), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[23][8]  (.Q (\o_values[23] [8] ), .CK (n_0_144), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[23][9]  (.Q (\o_values[23] [9] ), .CK (n_0_144), .D (sps__n37));
DFF_X1 \o_values_reg[23][10]  (.Q (\o_values[23] [10] ), .CK (n_0_144), .D (sps__n4));
DFF_X1 \o_values_reg[23][11]  (.Q (\o_values[23] [11] ), .CK (n_0_144), .D (sps__n10));
DFF_X1 \o_values_reg[23][12]  (.Q (\o_values[23] [12] ), .CK (n_0_144), .D (sps__n7));
DFF_X1 \o_values_reg[23][13]  (.Q (\o_values[23] [13] ), .CK (n_0_144), .D (sps__n1));
DFF_X1 \o_values_reg[23][14]  (.Q (\o_values[23] [14] ), .CK (n_0_144), .D (sps__n13));
DFF_X1 \o_values_reg[23][15]  (.Q (\o_values[23] [15] ), .CK (n_0_144), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[23]_reg  (.GCK (n_0_144), .CK (clk), .E (n_0_60), .SE (1'b0 ));
DFF_X1 \o_values_reg[24][0]  (.Q (\o_values[24] [0] ), .CK (n_0_143), .D (sps__n16));
DFF_X1 \o_values_reg[24][1]  (.Q (\o_values[24] [1] ), .CK (n_0_143), .D (sps__n25));
DFF_X1 \o_values_reg[24][2]  (.Q (\o_values[24] [2] ), .CK (n_0_143), .D (sps__n19));
DFF_X1 \o_values_reg[24][3]  (.Q (\o_values[24] [3] ), .CK (n_0_143), .D (sps__n28));
DFF_X1 \o_values_reg[24][4]  (.Q (\o_values[24] [4] ), .CK (n_0_143), .D (sps__n31));
DFF_X1 \o_values_reg[24][5]  (.Q (\o_values[24] [5] ), .CK (n_0_143), .D (sps__n34));
DFF_X1 \o_values_reg[24][6]  (.Q (\o_values[24] [6] ), .CK (n_0_143), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[24][7]  (.Q (\o_values[24] [7] ), .CK (n_0_143), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[24][8]  (.Q (\o_values[24] [8] ), .CK (n_0_143), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[24][9]  (.Q (\o_values[24] [9] ), .CK (n_0_143), .D (sps__n37));
DFF_X1 \o_values_reg[24][10]  (.Q (\o_values[24] [10] ), .CK (n_0_143), .D (sps__n4));
DFF_X1 \o_values_reg[24][11]  (.Q (\o_values[24] [11] ), .CK (n_0_143), .D (sps__n10));
DFF_X1 \o_values_reg[24][12]  (.Q (\o_values[24] [12] ), .CK (n_0_143), .D (sps__n7));
DFF_X1 \o_values_reg[24][13]  (.Q (\o_values[24] [13] ), .CK (n_0_143), .D (sps__n1));
DFF_X1 \o_values_reg[24][14]  (.Q (\o_values[24] [14] ), .CK (n_0_143), .D (sps__n13));
DFF_X1 \o_values_reg[24][15]  (.Q (\o_values[24] [15] ), .CK (n_0_143), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[24]_reg  (.GCK (n_0_143), .CK (clk), .E (n_0_59), .SE (1'b0 ));
DFF_X1 \o_values_reg[25][0]  (.Q (\o_values[25] [0] ), .CK (n_0_142), .D (sps__n16));
DFF_X1 \o_values_reg[25][1]  (.Q (\o_values[25] [1] ), .CK (n_0_142), .D (sps__n25));
DFF_X1 \o_values_reg[25][2]  (.Q (\o_values[25] [2] ), .CK (n_0_142), .D (sps__n19));
DFF_X1 \o_values_reg[25][3]  (.Q (\o_values[25] [3] ), .CK (n_0_142), .D (sps__n28));
DFF_X1 \o_values_reg[25][4]  (.Q (\o_values[25] [4] ), .CK (n_0_142), .D (sps__n31));
DFF_X1 \o_values_reg[25][5]  (.Q (\o_values[25] [5] ), .CK (n_0_142), .D (sps__n34));
DFF_X1 \o_values_reg[25][6]  (.Q (\o_values[25] [6] ), .CK (n_0_142), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[25][7]  (.Q (\o_values[25] [7] ), .CK (n_0_142), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[25][8]  (.Q (\o_values[25] [8] ), .CK (n_0_142), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[25][9]  (.Q (\o_values[25] [9] ), .CK (n_0_142), .D (sps__n37));
DFF_X1 \o_values_reg[25][10]  (.Q (\o_values[25] [10] ), .CK (n_0_142), .D (sps__n4));
DFF_X1 \o_values_reg[25][11]  (.Q (\o_values[25] [11] ), .CK (n_0_142), .D (sps__n10));
DFF_X1 \o_values_reg[25][12]  (.Q (\o_values[25] [12] ), .CK (n_0_142), .D (sps__n7));
DFF_X1 \o_values_reg[25][13]  (.Q (\o_values[25] [13] ), .CK (n_0_142), .D (sps__n1));
DFF_X1 \o_values_reg[25][14]  (.Q (\o_values[25] [14] ), .CK (n_0_142), .D (sps__n13));
DFF_X1 \o_values_reg[25][15]  (.Q (\o_values[25] [15] ), .CK (n_0_142), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[25]_reg  (.GCK (n_0_142), .CK (clk), .E (n_0_58), .SE (1'b0 ));
DFF_X1 \o_values_reg[26][0]  (.Q (\o_values[26] [0] ), .CK (n_0_141), .D (sps__n16));
DFF_X1 \o_values_reg[26][1]  (.Q (\o_values[26] [1] ), .CK (n_0_141), .D (sps__n25));
DFF_X1 \o_values_reg[26][2]  (.Q (\o_values[26] [2] ), .CK (n_0_141), .D (sps__n19));
DFF_X1 \o_values_reg[26][3]  (.Q (\o_values[26] [3] ), .CK (n_0_141), .D (sps__n28));
DFF_X1 \o_values_reg[26][4]  (.Q (\o_values[26] [4] ), .CK (n_0_141), .D (sps__n31));
DFF_X1 \o_values_reg[26][5]  (.Q (\o_values[26] [5] ), .CK (n_0_141), .D (sps__n34));
DFF_X1 \o_values_reg[26][6]  (.Q (\o_values[26] [6] ), .CK (n_0_141), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[26][7]  (.Q (\o_values[26] [7] ), .CK (n_0_141), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[26][8]  (.Q (\o_values[26] [8] ), .CK (n_0_141), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[26][9]  (.Q (\o_values[26] [9] ), .CK (n_0_141), .D (sps__n37));
DFF_X1 \o_values_reg[26][10]  (.Q (\o_values[26] [10] ), .CK (n_0_141), .D (sps__n4));
DFF_X1 \o_values_reg[26][11]  (.Q (\o_values[26] [11] ), .CK (n_0_141), .D (sps__n10));
DFF_X1 \o_values_reg[26][12]  (.Q (\o_values[26] [12] ), .CK (n_0_141), .D (sps__n7));
DFF_X1 \o_values_reg[26][13]  (.Q (\o_values[26] [13] ), .CK (n_0_141), .D (sps__n1));
DFF_X1 \o_values_reg[26][14]  (.Q (\o_values[26] [14] ), .CK (n_0_141), .D (sps__n13));
DFF_X1 \o_values_reg[26][15]  (.Q (\o_values[26] [15] ), .CK (n_0_141), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[26]_reg  (.GCK (n_0_141), .CK (clk), .E (n_0_57), .SE (1'b0 ));
DFF_X1 \o_values_reg[27][0]  (.Q (\o_values[27] [0] ), .CK (n_0_140), .D (sps__n16));
DFF_X1 \o_values_reg[27][1]  (.Q (\o_values[27] [1] ), .CK (n_0_140), .D (sps__n25));
DFF_X1 \o_values_reg[27][2]  (.Q (\o_values[27] [2] ), .CK (n_0_140), .D (sps__n19));
DFF_X1 \o_values_reg[27][3]  (.Q (\o_values[27] [3] ), .CK (n_0_140), .D (sps__n28));
DFF_X1 \o_values_reg[27][4]  (.Q (\o_values[27] [4] ), .CK (n_0_140), .D (sps__n31));
DFF_X1 \o_values_reg[27][5]  (.Q (\o_values[27] [5] ), .CK (n_0_140), .D (sps__n34));
DFF_X1 \o_values_reg[27][6]  (.Q (\o_values[27] [6] ), .CK (n_0_140), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[27][7]  (.Q (\o_values[27] [7] ), .CK (n_0_140), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[27][8]  (.Q (\o_values[27] [8] ), .CK (n_0_140), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[27][9]  (.Q (\o_values[27] [9] ), .CK (n_0_140), .D (sps__n37));
DFF_X1 \o_values_reg[27][10]  (.Q (\o_values[27] [10] ), .CK (n_0_140), .D (sps__n4));
DFF_X1 \o_values_reg[27][11]  (.Q (\o_values[27] [11] ), .CK (n_0_140), .D (sps__n10));
DFF_X1 \o_values_reg[27][12]  (.Q (\o_values[27] [12] ), .CK (n_0_140), .D (sps__n7));
DFF_X1 \o_values_reg[27][13]  (.Q (\o_values[27] [13] ), .CK (n_0_140), .D (sps__n1));
DFF_X1 \o_values_reg[27][14]  (.Q (\o_values[27] [14] ), .CK (n_0_140), .D (sps__n13));
DFF_X1 \o_values_reg[27][15]  (.Q (\o_values[27] [15] ), .CK (n_0_140), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[27]_reg  (.GCK (n_0_140), .CK (clk), .E (n_0_56), .SE (1'b0 ));
DFF_X1 \o_values_reg[28][0]  (.Q (\o_values[28] [0] ), .CK (n_0_139), .D (sps__n16));
DFF_X1 \o_values_reg[28][1]  (.Q (\o_values[28] [1] ), .CK (n_0_139), .D (sps__n25));
DFF_X1 \o_values_reg[28][2]  (.Q (\o_values[28] [2] ), .CK (n_0_139), .D (sps__n19));
DFF_X1 \o_values_reg[28][3]  (.Q (\o_values[28] [3] ), .CK (n_0_139), .D (sps__n28));
DFF_X1 \o_values_reg[28][4]  (.Q (\o_values[28] [4] ), .CK (n_0_139), .D (sps__n31));
DFF_X1 \o_values_reg[28][5]  (.Q (\o_values[28] [5] ), .CK (n_0_139), .D (sps__n34));
DFF_X1 \o_values_reg[28][6]  (.Q (\o_values[28] [6] ), .CK (n_0_139), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[28][7]  (.Q (\o_values[28] [7] ), .CK (n_0_139), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[28][8]  (.Q (\o_values[28] [8] ), .CK (n_0_139), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[28][9]  (.Q (\o_values[28] [9] ), .CK (n_0_139), .D (sps__n37));
DFF_X1 \o_values_reg[28][10]  (.Q (\o_values[28] [10] ), .CK (n_0_139), .D (sps__n4));
DFF_X1 \o_values_reg[28][11]  (.Q (\o_values[28] [11] ), .CK (n_0_139), .D (sps__n10));
DFF_X1 \o_values_reg[28][12]  (.Q (\o_values[28] [12] ), .CK (n_0_139), .D (sps__n7));
DFF_X1 \o_values_reg[28][13]  (.Q (\o_values[28] [13] ), .CK (n_0_139), .D (sps__n1));
DFF_X1 \o_values_reg[28][14]  (.Q (\o_values[28] [14] ), .CK (n_0_139), .D (sps__n13));
DFF_X1 \o_values_reg[28][15]  (.Q (\o_values[28] [15] ), .CK (n_0_139), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[28]_reg  (.GCK (n_0_139), .CK (clk), .E (n_0_55), .SE (1'b0 ));
DFF_X1 \o_values_reg[29][0]  (.Q (\o_values[29] [0] ), .CK (n_0_138), .D (sps__n16));
DFF_X1 \o_values_reg[29][1]  (.Q (\o_values[29] [1] ), .CK (n_0_138), .D (sps__n25));
DFF_X1 \o_values_reg[29][2]  (.Q (\o_values[29] [2] ), .CK (n_0_138), .D (sps__n19));
DFF_X1 \o_values_reg[29][3]  (.Q (\o_values[29] [3] ), .CK (n_0_138), .D (sps__n28));
DFF_X1 \o_values_reg[29][4]  (.Q (\o_values[29] [4] ), .CK (n_0_138), .D (sps__n31));
DFF_X1 \o_values_reg[29][5]  (.Q (\o_values[29] [5] ), .CK (n_0_138), .D (sps__n34));
DFF_X1 \o_values_reg[29][6]  (.Q (\o_values[29] [6] ), .CK (n_0_138), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[29][7]  (.Q (\o_values[29] [7] ), .CK (n_0_138), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[29][8]  (.Q (\o_values[29] [8] ), .CK (n_0_138), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[29][9]  (.Q (\o_values[29] [9] ), .CK (n_0_138), .D (sps__n37));
DFF_X1 \o_values_reg[29][10]  (.Q (\o_values[29] [10] ), .CK (n_0_138), .D (sps__n4));
DFF_X1 \o_values_reg[29][11]  (.Q (\o_values[29] [11] ), .CK (n_0_138), .D (sps__n10));
DFF_X1 \o_values_reg[29][12]  (.Q (\o_values[29] [12] ), .CK (n_0_138), .D (sps__n7));
DFF_X1 \o_values_reg[29][13]  (.Q (\o_values[29] [13] ), .CK (n_0_138), .D (sps__n1));
DFF_X1 \o_values_reg[29][14]  (.Q (\o_values[29] [14] ), .CK (n_0_138), .D (sps__n13));
DFF_X1 \o_values_reg[29][15]  (.Q (\o_values[29] [15] ), .CK (n_0_138), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[29]_reg  (.GCK (n_0_138), .CK (clk), .E (n_0_54), .SE (1'b0 ));
DFF_X1 \o_values_reg[30][0]  (.Q (\o_values[30] [0] ), .CK (n_0_137), .D (sps__n16));
DFF_X1 \o_values_reg[30][1]  (.Q (\o_values[30] [1] ), .CK (n_0_137), .D (sps__n25));
DFF_X1 \o_values_reg[30][2]  (.Q (\o_values[30] [2] ), .CK (n_0_137), .D (sps__n19));
DFF_X1 \o_values_reg[30][3]  (.Q (\o_values[30] [3] ), .CK (n_0_137), .D (sps__n28));
DFF_X1 \o_values_reg[30][4]  (.Q (\o_values[30] [4] ), .CK (n_0_137), .D (sps__n31));
DFF_X1 \o_values_reg[30][5]  (.Q (\o_values[30] [5] ), .CK (n_0_137), .D (sps__n34));
DFF_X1 \o_values_reg[30][6]  (.Q (\o_values[30] [6] ), .CK (n_0_137), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[30][7]  (.Q (\o_values[30] [7] ), .CK (n_0_137), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[30][8]  (.Q (\o_values[30] [8] ), .CK (n_0_137), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[30][9]  (.Q (\o_values[30] [9] ), .CK (n_0_137), .D (sps__n37));
DFF_X1 \o_values_reg[30][10]  (.Q (\o_values[30] [10] ), .CK (n_0_137), .D (sps__n4));
DFF_X1 \o_values_reg[30][11]  (.Q (\o_values[30] [11] ), .CK (n_0_137), .D (sps__n10));
DFF_X1 \o_values_reg[30][12]  (.Q (\o_values[30] [12] ), .CK (n_0_137), .D (sps__n7));
DFF_X1 \o_values_reg[30][13]  (.Q (\o_values[30] [13] ), .CK (n_0_137), .D (sps__n1));
DFF_X1 \o_values_reg[30][14]  (.Q (\o_values[30] [14] ), .CK (n_0_137), .D (sps__n13));
DFF_X1 \o_values_reg[30][15]  (.Q (\o_values[30] [15] ), .CK (n_0_137), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[30]_reg  (.GCK (n_0_137), .CK (clk), .E (n_0_53), .SE (1'b0 ));
DFF_X1 \o_values_reg[31][0]  (.Q (\o_values[31] [0] ), .CK (n_0_136), .D (sps__n16));
DFF_X1 \o_values_reg[31][1]  (.Q (\o_values[31] [1] ), .CK (n_0_136), .D (sps__n25));
DFF_X1 \o_values_reg[31][2]  (.Q (\o_values[31] [2] ), .CK (n_0_136), .D (sps__n19));
DFF_X1 \o_values_reg[31][3]  (.Q (\o_values[31] [3] ), .CK (n_0_136), .D (sps__n28));
DFF_X1 \o_values_reg[31][4]  (.Q (\o_values[31] [4] ), .CK (n_0_136), .D (sps__n31));
DFF_X1 \o_values_reg[31][5]  (.Q (\o_values[31] [5] ), .CK (n_0_136), .D (sps__n34));
DFF_X1 \o_values_reg[31][6]  (.Q (\o_values[31] [6] ), .CK (n_0_136), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[31][7]  (.Q (\o_values[31] [7] ), .CK (n_0_136), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[31][8]  (.Q (\o_values[31] [8] ), .CK (n_0_136), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[31][9]  (.Q (\o_values[31] [9] ), .CK (n_0_136), .D (sps__n37));
DFF_X1 \o_values_reg[31][10]  (.Q (\o_values[31] [10] ), .CK (n_0_136), .D (sps__n4));
DFF_X1 \o_values_reg[31][11]  (.Q (\o_values[31] [11] ), .CK (n_0_136), .D (sps__n10));
DFF_X1 \o_values_reg[31][12]  (.Q (\o_values[31] [12] ), .CK (n_0_136), .D (sps__n7));
DFF_X1 \o_values_reg[31][13]  (.Q (\o_values[31] [13] ), .CK (n_0_136), .D (sps__n1));
DFF_X1 \o_values_reg[31][14]  (.Q (\o_values[31] [14] ), .CK (n_0_136), .D (sps__n13));
DFF_X1 \o_values_reg[31][15]  (.Q (\o_values[31] [15] ), .CK (n_0_136), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[31]_reg  (.GCK (n_0_136), .CK (clk), .E (n_0_52), .SE (1'b0 ));
DFF_X1 \o_values_reg[32][0]  (.Q (\o_values[32] [0] ), .CK (n_0_135), .D (sps__n16));
DFF_X1 \o_values_reg[32][1]  (.Q (\o_values[32] [1] ), .CK (n_0_135), .D (sps__n25));
DFF_X1 \o_values_reg[32][2]  (.Q (\o_values[32] [2] ), .CK (n_0_135), .D (sps__n19));
DFF_X1 \o_values_reg[32][3]  (.Q (\o_values[32] [3] ), .CK (n_0_135), .D (sps__n28));
DFF_X1 \o_values_reg[32][4]  (.Q (\o_values[32] [4] ), .CK (n_0_135), .D (sps__n31));
DFF_X1 \o_values_reg[32][5]  (.Q (\o_values[32] [5] ), .CK (n_0_135), .D (sps__n34));
DFF_X1 \o_values_reg[32][6]  (.Q (\o_values[32] [6] ), .CK (n_0_135), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[32][7]  (.Q (\o_values[32] [7] ), .CK (n_0_135), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[32][8]  (.Q (\o_values[32] [8] ), .CK (n_0_135), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[32][9]  (.Q (\o_values[32] [9] ), .CK (n_0_135), .D (sps__n37));
DFF_X1 \o_values_reg[32][10]  (.Q (\o_values[32] [10] ), .CK (n_0_135), .D (sps__n4));
DFF_X1 \o_values_reg[32][11]  (.Q (\o_values[32] [11] ), .CK (n_0_135), .D (sps__n10));
DFF_X1 \o_values_reg[32][12]  (.Q (\o_values[32] [12] ), .CK (n_0_135), .D (sps__n7));
DFF_X1 \o_values_reg[32][13]  (.Q (\o_values[32] [13] ), .CK (n_0_135), .D (sps__n1));
DFF_X1 \o_values_reg[32][14]  (.Q (\o_values[32] [14] ), .CK (n_0_135), .D (sps__n13));
DFF_X1 \o_values_reg[32][15]  (.Q (\o_values[32] [15] ), .CK (n_0_135), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[32]_reg  (.GCK (n_0_135), .CK (clk), .E (n_0_51), .SE (1'b0 ));
DFF_X1 \o_values_reg[33][0]  (.Q (\o_values[33] [0] ), .CK (n_0_134), .D (sps__n16));
DFF_X1 \o_values_reg[33][1]  (.Q (\o_values[33] [1] ), .CK (n_0_134), .D (sps__n25));
DFF_X1 \o_values_reg[33][2]  (.Q (\o_values[33] [2] ), .CK (n_0_134), .D (sps__n19));
DFF_X1 \o_values_reg[33][3]  (.Q (\o_values[33] [3] ), .CK (n_0_134), .D (sps__n28));
DFF_X1 \o_values_reg[33][4]  (.Q (\o_values[33] [4] ), .CK (n_0_134), .D (sps__n31));
DFF_X1 \o_values_reg[33][5]  (.Q (\o_values[33] [5] ), .CK (n_0_134), .D (sps__n34));
DFF_X1 \o_values_reg[33][6]  (.Q (\o_values[33] [6] ), .CK (n_0_134), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[33][7]  (.Q (\o_values[33] [7] ), .CK (n_0_134), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[33][8]  (.Q (\o_values[33] [8] ), .CK (n_0_134), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[33][9]  (.Q (\o_values[33] [9] ), .CK (n_0_134), .D (sps__n37));
DFF_X1 \o_values_reg[33][10]  (.Q (\o_values[33] [10] ), .CK (n_0_134), .D (sps__n4));
DFF_X1 \o_values_reg[33][11]  (.Q (\o_values[33] [11] ), .CK (n_0_134), .D (sps__n10));
DFF_X1 \o_values_reg[33][12]  (.Q (\o_values[33] [12] ), .CK (n_0_134), .D (sps__n7));
DFF_X1 \o_values_reg[33][13]  (.Q (\o_values[33] [13] ), .CK (n_0_134), .D (sps__n1));
DFF_X1 \o_values_reg[33][14]  (.Q (\o_values[33] [14] ), .CK (n_0_134), .D (sps__n13));
DFF_X1 \o_values_reg[33][15]  (.Q (\o_values[33] [15] ), .CK (n_0_134), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[33]_reg  (.GCK (n_0_134), .CK (clk), .E (n_0_50), .SE (1'b0 ));
DFF_X1 \o_values_reg[34][0]  (.Q (\o_values[34] [0] ), .CK (n_0_133), .D (sps__n16));
DFF_X1 \o_values_reg[34][1]  (.Q (\o_values[34] [1] ), .CK (n_0_133), .D (sps__n25));
DFF_X1 \o_values_reg[34][2]  (.Q (\o_values[34] [2] ), .CK (n_0_133), .D (sps__n19));
DFF_X1 \o_values_reg[34][3]  (.Q (\o_values[34] [3] ), .CK (n_0_133), .D (sps__n28));
DFF_X1 \o_values_reg[34][4]  (.Q (\o_values[34] [4] ), .CK (n_0_133), .D (sps__n31));
DFF_X1 \o_values_reg[34][5]  (.Q (\o_values[34] [5] ), .CK (n_0_133), .D (sps__n34));
DFF_X1 \o_values_reg[34][6]  (.Q (\o_values[34] [6] ), .CK (n_0_133), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[34][7]  (.Q (\o_values[34] [7] ), .CK (n_0_133), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[34][8]  (.Q (\o_values[34] [8] ), .CK (n_0_133), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[34][9]  (.Q (\o_values[34] [9] ), .CK (n_0_133), .D (sps__n37));
DFF_X1 \o_values_reg[34][10]  (.Q (\o_values[34] [10] ), .CK (n_0_133), .D (sps__n4));
DFF_X1 \o_values_reg[34][11]  (.Q (\o_values[34] [11] ), .CK (n_0_133), .D (sps__n10));
DFF_X1 \o_values_reg[34][12]  (.Q (\o_values[34] [12] ), .CK (n_0_133), .D (sps__n7));
DFF_X1 \o_values_reg[34][13]  (.Q (\o_values[34] [13] ), .CK (n_0_133), .D (sps__n1));
DFF_X1 \o_values_reg[34][14]  (.Q (\o_values[34] [14] ), .CK (n_0_133), .D (sps__n13));
DFF_X1 \o_values_reg[34][15]  (.Q (\o_values[34] [15] ), .CK (n_0_133), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[34]_reg  (.GCK (n_0_133), .CK (clk), .E (n_0_49), .SE (1'b0 ));
DFF_X1 \o_values_reg[35][0]  (.Q (\o_values[35] [0] ), .CK (n_0_132), .D (sps__n16));
DFF_X1 \o_values_reg[35][1]  (.Q (\o_values[35] [1] ), .CK (n_0_132), .D (sps__n25));
DFF_X1 \o_values_reg[35][2]  (.Q (\o_values[35] [2] ), .CK (n_0_132), .D (sps__n19));
DFF_X1 \o_values_reg[35][3]  (.Q (\o_values[35] [3] ), .CK (n_0_132), .D (sps__n28));
DFF_X1 \o_values_reg[35][4]  (.Q (\o_values[35] [4] ), .CK (n_0_132), .D (sps__n31));
DFF_X1 \o_values_reg[35][5]  (.Q (\o_values[35] [5] ), .CK (n_0_132), .D (sps__n34));
DFF_X1 \o_values_reg[35][6]  (.Q (\o_values[35] [6] ), .CK (n_0_132), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[35][7]  (.Q (\o_values[35] [7] ), .CK (n_0_132), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[35][8]  (.Q (\o_values[35] [8] ), .CK (n_0_132), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[35][9]  (.Q (\o_values[35] [9] ), .CK (n_0_132), .D (sps__n37));
DFF_X1 \o_values_reg[35][10]  (.Q (\o_values[35] [10] ), .CK (n_0_132), .D (sps__n4));
DFF_X1 \o_values_reg[35][11]  (.Q (\o_values[35] [11] ), .CK (n_0_132), .D (sps__n10));
DFF_X1 \o_values_reg[35][12]  (.Q (\o_values[35] [12] ), .CK (n_0_132), .D (sps__n7));
DFF_X1 \o_values_reg[35][13]  (.Q (\o_values[35] [13] ), .CK (n_0_132), .D (sps__n1));
DFF_X1 \o_values_reg[35][14]  (.Q (\o_values[35] [14] ), .CK (n_0_132), .D (sps__n13));
DFF_X1 \o_values_reg[35][15]  (.Q (\o_values[35] [15] ), .CK (n_0_132), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[35]_reg  (.GCK (n_0_132), .CK (clk), .E (n_0_48), .SE (1'b0 ));
DFF_X1 \o_values_reg[36][0]  (.Q (\o_values[36] [0] ), .CK (n_0_131), .D (sps__n16));
DFF_X1 \o_values_reg[36][1]  (.Q (\o_values[36] [1] ), .CK (n_0_131), .D (sps__n25));
DFF_X1 \o_values_reg[36][2]  (.Q (\o_values[36] [2] ), .CK (n_0_131), .D (sps__n19));
DFF_X1 \o_values_reg[36][3]  (.Q (\o_values[36] [3] ), .CK (n_0_131), .D (sps__n28));
DFF_X1 \o_values_reg[36][4]  (.Q (\o_values[36] [4] ), .CK (n_0_131), .D (sps__n31));
DFF_X1 \o_values_reg[36][5]  (.Q (\o_values[36] [5] ), .CK (n_0_131), .D (sps__n34));
DFF_X1 \o_values_reg[36][6]  (.Q (\o_values[36] [6] ), .CK (n_0_131), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[36][7]  (.Q (\o_values[36] [7] ), .CK (n_0_131), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[36][8]  (.Q (\o_values[36] [8] ), .CK (n_0_131), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[36][9]  (.Q (\o_values[36] [9] ), .CK (n_0_131), .D (sps__n37));
DFF_X1 \o_values_reg[36][10]  (.Q (\o_values[36] [10] ), .CK (n_0_131), .D (sps__n4));
DFF_X1 \o_values_reg[36][11]  (.Q (\o_values[36] [11] ), .CK (n_0_131), .D (sps__n10));
DFF_X1 \o_values_reg[36][12]  (.Q (\o_values[36] [12] ), .CK (n_0_131), .D (sps__n7));
DFF_X1 \o_values_reg[36][13]  (.Q (\o_values[36] [13] ), .CK (n_0_131), .D (sps__n1));
DFF_X1 \o_values_reg[36][14]  (.Q (\o_values[36] [14] ), .CK (n_0_131), .D (sps__n13));
DFF_X1 \o_values_reg[36][15]  (.Q (\o_values[36] [15] ), .CK (n_0_131), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[36]_reg  (.GCK (n_0_131), .CK (clk), .E (n_0_47), .SE (1'b0 ));
DFF_X1 \o_values_reg[37][0]  (.Q (\o_values[37] [0] ), .CK (n_0_130), .D (sps__n16));
DFF_X1 \o_values_reg[37][1]  (.Q (\o_values[37] [1] ), .CK (n_0_130), .D (sps__n25));
DFF_X1 \o_values_reg[37][2]  (.Q (\o_values[37] [2] ), .CK (n_0_130), .D (sps__n19));
DFF_X1 \o_values_reg[37][3]  (.Q (\o_values[37] [3] ), .CK (n_0_130), .D (sps__n28));
DFF_X1 \o_values_reg[37][4]  (.Q (\o_values[37] [4] ), .CK (n_0_130), .D (sps__n31));
DFF_X1 \o_values_reg[37][5]  (.Q (\o_values[37] [5] ), .CK (n_0_130), .D (sps__n34));
DFF_X1 \o_values_reg[37][6]  (.Q (\o_values[37] [6] ), .CK (n_0_130), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[37][7]  (.Q (\o_values[37] [7] ), .CK (n_0_130), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[37][8]  (.Q (\o_values[37] [8] ), .CK (n_0_130), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[37][9]  (.Q (\o_values[37] [9] ), .CK (n_0_130), .D (sps__n37));
DFF_X1 \o_values_reg[37][10]  (.Q (\o_values[37] [10] ), .CK (n_0_130), .D (sps__n4));
DFF_X1 \o_values_reg[37][11]  (.Q (\o_values[37] [11] ), .CK (n_0_130), .D (sps__n10));
DFF_X1 \o_values_reg[37][12]  (.Q (\o_values[37] [12] ), .CK (n_0_130), .D (sps__n7));
DFF_X1 \o_values_reg[37][13]  (.Q (\o_values[37] [13] ), .CK (n_0_130), .D (sps__n1));
DFF_X1 \o_values_reg[37][14]  (.Q (\o_values[37] [14] ), .CK (n_0_130), .D (sps__n13));
DFF_X1 \o_values_reg[37][15]  (.Q (\o_values[37] [15] ), .CK (n_0_130), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[37]_reg  (.GCK (n_0_130), .CK (clk), .E (n_0_46), .SE (1'b0 ));
DFF_X1 \o_values_reg[38][0]  (.Q (\o_values[38] [0] ), .CK (n_0_129), .D (sps__n16));
DFF_X1 \o_values_reg[38][1]  (.Q (\o_values[38] [1] ), .CK (n_0_129), .D (sps__n25));
DFF_X1 \o_values_reg[38][2]  (.Q (\o_values[38] [2] ), .CK (n_0_129), .D (sps__n19));
DFF_X1 \o_values_reg[38][3]  (.Q (\o_values[38] [3] ), .CK (n_0_129), .D (sps__n28));
DFF_X1 \o_values_reg[38][4]  (.Q (\o_values[38] [4] ), .CK (n_0_129), .D (sps__n31));
DFF_X1 \o_values_reg[38][5]  (.Q (\o_values[38] [5] ), .CK (n_0_129), .D (sps__n34));
DFF_X1 \o_values_reg[38][6]  (.Q (\o_values[38] [6] ), .CK (n_0_129), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[38][7]  (.Q (\o_values[38] [7] ), .CK (n_0_129), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[38][8]  (.Q (\o_values[38] [8] ), .CK (n_0_129), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[38][9]  (.Q (\o_values[38] [9] ), .CK (n_0_129), .D (sps__n37));
DFF_X1 \o_values_reg[38][10]  (.Q (\o_values[38] [10] ), .CK (n_0_129), .D (sps__n4));
DFF_X1 \o_values_reg[38][11]  (.Q (\o_values[38] [11] ), .CK (n_0_129), .D (sps__n10));
DFF_X1 \o_values_reg[38][12]  (.Q (\o_values[38] [12] ), .CK (n_0_129), .D (sps__n7));
DFF_X1 \o_values_reg[38][13]  (.Q (\o_values[38] [13] ), .CK (n_0_129), .D (sps__n1));
DFF_X1 \o_values_reg[38][14]  (.Q (\o_values[38] [14] ), .CK (n_0_129), .D (sps__n13));
DFF_X1 \o_values_reg[38][15]  (.Q (\o_values[38] [15] ), .CK (n_0_129), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[38]_reg  (.GCK (n_0_129), .CK (clk), .E (n_0_45), .SE (1'b0 ));
DFF_X1 \o_values_reg[39][0]  (.Q (\o_values[39] [0] ), .CK (n_0_128), .D (sps__n16));
DFF_X1 \o_values_reg[39][1]  (.Q (\o_values[39] [1] ), .CK (n_0_128), .D (sps__n25));
DFF_X1 \o_values_reg[39][2]  (.Q (\o_values[39] [2] ), .CK (n_0_128), .D (sps__n19));
DFF_X1 \o_values_reg[39][3]  (.Q (\o_values[39] [3] ), .CK (n_0_128), .D (sps__n28));
DFF_X1 \o_values_reg[39][4]  (.Q (\o_values[39] [4] ), .CK (n_0_128), .D (sps__n31));
DFF_X1 \o_values_reg[39][5]  (.Q (\o_values[39] [5] ), .CK (n_0_128), .D (sps__n34));
DFF_X1 \o_values_reg[39][6]  (.Q (\o_values[39] [6] ), .CK (n_0_128), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[39][7]  (.Q (\o_values[39] [7] ), .CK (n_0_128), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[39][8]  (.Q (\o_values[39] [8] ), .CK (n_0_128), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[39][9]  (.Q (\o_values[39] [9] ), .CK (n_0_128), .D (sps__n37));
DFF_X1 \o_values_reg[39][10]  (.Q (\o_values[39] [10] ), .CK (n_0_128), .D (sps__n4));
DFF_X1 \o_values_reg[39][11]  (.Q (\o_values[39] [11] ), .CK (n_0_128), .D (sps__n10));
DFF_X1 \o_values_reg[39][12]  (.Q (\o_values[39] [12] ), .CK (n_0_128), .D (sps__n7));
DFF_X1 \o_values_reg[39][13]  (.Q (\o_values[39] [13] ), .CK (n_0_128), .D (sps__n1));
DFF_X1 \o_values_reg[39][14]  (.Q (\o_values[39] [14] ), .CK (n_0_128), .D (sps__n13));
DFF_X1 \o_values_reg[39][15]  (.Q (\o_values[39] [15] ), .CK (n_0_128), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[39]_reg  (.GCK (n_0_128), .CK (clk), .E (n_0_44), .SE (1'b0 ));
DFF_X1 \o_values_reg[40][0]  (.Q (\o_values[40] [0] ), .CK (n_0_127), .D (sps__n16));
DFF_X1 \o_values_reg[40][1]  (.Q (\o_values[40] [1] ), .CK (n_0_127), .D (sps__n25));
DFF_X1 \o_values_reg[40][2]  (.Q (\o_values[40] [2] ), .CK (n_0_127), .D (sps__n19));
DFF_X1 \o_values_reg[40][3]  (.Q (\o_values[40] [3] ), .CK (n_0_127), .D (sps__n28));
DFF_X1 \o_values_reg[40][4]  (.Q (\o_values[40] [4] ), .CK (n_0_127), .D (sps__n31));
DFF_X1 \o_values_reg[40][5]  (.Q (\o_values[40] [5] ), .CK (n_0_127), .D (sps__n34));
DFF_X1 \o_values_reg[40][6]  (.Q (\o_values[40] [6] ), .CK (n_0_127), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[40][7]  (.Q (\o_values[40] [7] ), .CK (n_0_127), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[40][8]  (.Q (\o_values[40] [8] ), .CK (n_0_127), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[40][9]  (.Q (\o_values[40] [9] ), .CK (n_0_127), .D (sps__n37));
DFF_X1 \o_values_reg[40][10]  (.Q (\o_values[40] [10] ), .CK (n_0_127), .D (sps__n4));
DFF_X1 \o_values_reg[40][11]  (.Q (\o_values[40] [11] ), .CK (n_0_127), .D (sps__n10));
DFF_X1 \o_values_reg[40][12]  (.Q (\o_values[40] [12] ), .CK (n_0_127), .D (sps__n7));
DFF_X1 \o_values_reg[40][13]  (.Q (\o_values[40] [13] ), .CK (n_0_127), .D (sps__n1));
DFF_X1 \o_values_reg[40][14]  (.Q (\o_values[40] [14] ), .CK (n_0_127), .D (sps__n13));
DFF_X1 \o_values_reg[40][15]  (.Q (\o_values[40] [15] ), .CK (n_0_127), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[40]_reg  (.GCK (n_0_127), .CK (clk), .E (n_0_43), .SE (1'b0 ));
DFF_X1 \o_values_reg[41][0]  (.Q (\o_values[41] [0] ), .CK (n_0_126), .D (sps__n16));
DFF_X1 \o_values_reg[41][1]  (.Q (\o_values[41] [1] ), .CK (n_0_126), .D (sps__n25));
DFF_X1 \o_values_reg[41][2]  (.Q (\o_values[41] [2] ), .CK (n_0_126), .D (sps__n19));
DFF_X1 \o_values_reg[41][3]  (.Q (\o_values[41] [3] ), .CK (n_0_126), .D (sps__n28));
DFF_X1 \o_values_reg[41][4]  (.Q (\o_values[41] [4] ), .CK (n_0_126), .D (sps__n31));
DFF_X1 \o_values_reg[41][5]  (.Q (\o_values[41] [5] ), .CK (n_0_126), .D (sps__n34));
DFF_X1 \o_values_reg[41][6]  (.Q (\o_values[41] [6] ), .CK (n_0_126), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[41][7]  (.Q (\o_values[41] [7] ), .CK (n_0_126), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[41][8]  (.Q (\o_values[41] [8] ), .CK (n_0_126), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[41][9]  (.Q (\o_values[41] [9] ), .CK (n_0_126), .D (sps__n37));
DFF_X1 \o_values_reg[41][10]  (.Q (\o_values[41] [10] ), .CK (n_0_126), .D (sps__n4));
DFF_X1 \o_values_reg[41][11]  (.Q (\o_values[41] [11] ), .CK (n_0_126), .D (sps__n10));
DFF_X1 \o_values_reg[41][12]  (.Q (\o_values[41] [12] ), .CK (n_0_126), .D (sps__n7));
DFF_X1 \o_values_reg[41][13]  (.Q (\o_values[41] [13] ), .CK (n_0_126), .D (sps__n1));
DFF_X1 \o_values_reg[41][14]  (.Q (\o_values[41] [14] ), .CK (n_0_126), .D (sps__n13));
DFF_X1 \o_values_reg[41][15]  (.Q (\o_values[41] [15] ), .CK (n_0_126), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[41]_reg  (.GCK (n_0_126), .CK (clk), .E (n_0_42), .SE (1'b0 ));
DFF_X1 \o_values_reg[42][0]  (.Q (\o_values[42] [0] ), .CK (n_0_125), .D (sps__n16));
DFF_X1 \o_values_reg[42][1]  (.Q (\o_values[42] [1] ), .CK (n_0_125), .D (sps__n25));
DFF_X1 \o_values_reg[42][2]  (.Q (\o_values[42] [2] ), .CK (n_0_125), .D (sps__n19));
DFF_X1 \o_values_reg[42][3]  (.Q (\o_values[42] [3] ), .CK (n_0_125), .D (sps__n28));
DFF_X1 \o_values_reg[42][4]  (.Q (\o_values[42] [4] ), .CK (n_0_125), .D (sps__n31));
DFF_X1 \o_values_reg[42][5]  (.Q (\o_values[42] [5] ), .CK (n_0_125), .D (sps__n34));
DFF_X1 \o_values_reg[42][6]  (.Q (\o_values[42] [6] ), .CK (n_0_125), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[42][7]  (.Q (\o_values[42] [7] ), .CK (n_0_125), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[42][8]  (.Q (\o_values[42] [8] ), .CK (n_0_125), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[42][9]  (.Q (\o_values[42] [9] ), .CK (n_0_125), .D (sps__n37));
DFF_X1 \o_values_reg[42][10]  (.Q (\o_values[42] [10] ), .CK (n_0_125), .D (sps__n4));
DFF_X1 \o_values_reg[42][11]  (.Q (\o_values[42] [11] ), .CK (n_0_125), .D (sps__n10));
DFF_X1 \o_values_reg[42][12]  (.Q (\o_values[42] [12] ), .CK (n_0_125), .D (sps__n7));
DFF_X1 \o_values_reg[42][13]  (.Q (\o_values[42] [13] ), .CK (n_0_125), .D (sps__n1));
DFF_X1 \o_values_reg[42][14]  (.Q (\o_values[42] [14] ), .CK (n_0_125), .D (sps__n13));
DFF_X1 \o_values_reg[42][15]  (.Q (\o_values[42] [15] ), .CK (n_0_125), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[42]_reg  (.GCK (n_0_125), .CK (clk), .E (n_0_41), .SE (1'b0 ));
DFF_X1 \o_values_reg[43][0]  (.Q (\o_values[43] [0] ), .CK (n_0_124), .D (sps__n16));
DFF_X1 \o_values_reg[43][1]  (.Q (\o_values[43] [1] ), .CK (n_0_124), .D (sps__n25));
DFF_X1 \o_values_reg[43][2]  (.Q (\o_values[43] [2] ), .CK (n_0_124), .D (sps__n19));
DFF_X1 \o_values_reg[43][3]  (.Q (\o_values[43] [3] ), .CK (n_0_124), .D (sps__n28));
DFF_X1 \o_values_reg[43][4]  (.Q (\o_values[43] [4] ), .CK (n_0_124), .D (sps__n31));
DFF_X1 \o_values_reg[43][5]  (.Q (\o_values[43] [5] ), .CK (n_0_124), .D (sps__n34));
DFF_X1 \o_values_reg[43][6]  (.Q (\o_values[43] [6] ), .CK (n_0_124), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[43][7]  (.Q (\o_values[43] [7] ), .CK (n_0_124), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[43][8]  (.Q (\o_values[43] [8] ), .CK (n_0_124), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[43][9]  (.Q (\o_values[43] [9] ), .CK (n_0_124), .D (sps__n37));
DFF_X1 \o_values_reg[43][10]  (.Q (\o_values[43] [10] ), .CK (n_0_124), .D (sps__n4));
DFF_X1 \o_values_reg[43][11]  (.Q (\o_values[43] [11] ), .CK (n_0_124), .D (sps__n10));
DFF_X1 \o_values_reg[43][12]  (.Q (\o_values[43] [12] ), .CK (n_0_124), .D (sps__n7));
DFF_X1 \o_values_reg[43][13]  (.Q (\o_values[43] [13] ), .CK (n_0_124), .D (sps__n1));
DFF_X1 \o_values_reg[43][14]  (.Q (\o_values[43] [14] ), .CK (n_0_124), .D (sps__n13));
DFF_X1 \o_values_reg[43][15]  (.Q (\o_values[43] [15] ), .CK (n_0_124), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[43]_reg  (.GCK (n_0_124), .CK (clk), .E (n_0_40), .SE (1'b0 ));
DFF_X1 \o_values_reg[44][0]  (.Q (\o_values[44] [0] ), .CK (n_0_123), .D (sps__n16));
DFF_X1 \o_values_reg[44][1]  (.Q (\o_values[44] [1] ), .CK (n_0_123), .D (sps__n25));
DFF_X1 \o_values_reg[44][2]  (.Q (\o_values[44] [2] ), .CK (n_0_123), .D (sps__n19));
DFF_X1 \o_values_reg[44][3]  (.Q (\o_values[44] [3] ), .CK (n_0_123), .D (sps__n28));
DFF_X1 \o_values_reg[44][4]  (.Q (\o_values[44] [4] ), .CK (n_0_123), .D (sps__n31));
DFF_X1 \o_values_reg[44][5]  (.Q (\o_values[44] [5] ), .CK (n_0_123), .D (sps__n34));
DFF_X1 \o_values_reg[44][6]  (.Q (\o_values[44] [6] ), .CK (n_0_123), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[44][7]  (.Q (\o_values[44] [7] ), .CK (n_0_123), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[44][8]  (.Q (\o_values[44] [8] ), .CK (n_0_123), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[44][9]  (.Q (\o_values[44] [9] ), .CK (n_0_123), .D (sps__n37));
DFF_X1 \o_values_reg[44][10]  (.Q (\o_values[44] [10] ), .CK (n_0_123), .D (sps__n4));
DFF_X1 \o_values_reg[44][11]  (.Q (\o_values[44] [11] ), .CK (n_0_123), .D (sps__n10));
DFF_X1 \o_values_reg[44][12]  (.Q (\o_values[44] [12] ), .CK (n_0_123), .D (sps__n7));
DFF_X1 \o_values_reg[44][13]  (.Q (\o_values[44] [13] ), .CK (n_0_123), .D (sps__n1));
DFF_X1 \o_values_reg[44][14]  (.Q (\o_values[44] [14] ), .CK (n_0_123), .D (sps__n13));
DFF_X1 \o_values_reg[44][15]  (.Q (\o_values[44] [15] ), .CK (n_0_123), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[44]_reg  (.GCK (n_0_123), .CK (clk), .E (n_0_39), .SE (1'b0 ));
DFF_X1 \o_values_reg[45][0]  (.Q (\o_values[45] [0] ), .CK (n_0_122), .D (sps__n16));
DFF_X1 \o_values_reg[45][1]  (.Q (\o_values[45] [1] ), .CK (n_0_122), .D (sps__n25));
DFF_X1 \o_values_reg[45][2]  (.Q (\o_values[45] [2] ), .CK (n_0_122), .D (sps__n19));
DFF_X1 \o_values_reg[45][3]  (.Q (\o_values[45] [3] ), .CK (n_0_122), .D (sps__n28));
DFF_X1 \o_values_reg[45][4]  (.Q (\o_values[45] [4] ), .CK (n_0_122), .D (sps__n31));
DFF_X1 \o_values_reg[45][5]  (.Q (\o_values[45] [5] ), .CK (n_0_122), .D (sps__n34));
DFF_X1 \o_values_reg[45][6]  (.Q (\o_values[45] [6] ), .CK (n_0_122), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[45][7]  (.Q (\o_values[45] [7] ), .CK (n_0_122), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[45][8]  (.Q (\o_values[45] [8] ), .CK (n_0_122), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[45][9]  (.Q (\o_values[45] [9] ), .CK (n_0_122), .D (sps__n37));
DFF_X1 \o_values_reg[45][10]  (.Q (\o_values[45] [10] ), .CK (n_0_122), .D (sps__n4));
DFF_X1 \o_values_reg[45][11]  (.Q (\o_values[45] [11] ), .CK (n_0_122), .D (sps__n10));
DFF_X1 \o_values_reg[45][12]  (.Q (\o_values[45] [12] ), .CK (n_0_122), .D (sps__n7));
DFF_X1 \o_values_reg[45][13]  (.Q (\o_values[45] [13] ), .CK (n_0_122), .D (sps__n1));
DFF_X1 \o_values_reg[45][14]  (.Q (\o_values[45] [14] ), .CK (n_0_122), .D (sps__n13));
DFF_X1 \o_values_reg[45][15]  (.Q (\o_values[45] [15] ), .CK (n_0_122), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[45]_reg  (.GCK (n_0_122), .CK (clk), .E (n_0_38), .SE (1'b0 ));
DFF_X1 \o_values_reg[46][0]  (.Q (\o_values[46] [0] ), .CK (n_0_121), .D (sps__n16));
DFF_X1 \o_values_reg[46][1]  (.Q (\o_values[46] [1] ), .CK (n_0_121), .D (sps__n25));
DFF_X1 \o_values_reg[46][2]  (.Q (\o_values[46] [2] ), .CK (n_0_121), .D (sps__n19));
DFF_X1 \o_values_reg[46][3]  (.Q (\o_values[46] [3] ), .CK (n_0_121), .D (sps__n28));
DFF_X1 \o_values_reg[46][4]  (.Q (\o_values[46] [4] ), .CK (n_0_121), .D (sps__n31));
DFF_X1 \o_values_reg[46][5]  (.Q (\o_values[46] [5] ), .CK (n_0_121), .D (sps__n34));
DFF_X1 \o_values_reg[46][6]  (.Q (\o_values[46] [6] ), .CK (n_0_121), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[46][7]  (.Q (\o_values[46] [7] ), .CK (n_0_121), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[46][8]  (.Q (\o_values[46] [8] ), .CK (n_0_121), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[46][9]  (.Q (\o_values[46] [9] ), .CK (n_0_121), .D (sps__n37));
DFF_X1 \o_values_reg[46][10]  (.Q (\o_values[46] [10] ), .CK (n_0_121), .D (sps__n4));
DFF_X1 \o_values_reg[46][11]  (.Q (\o_values[46] [11] ), .CK (n_0_121), .D (sps__n10));
DFF_X1 \o_values_reg[46][12]  (.Q (\o_values[46] [12] ), .CK (n_0_121), .D (sps__n7));
DFF_X1 \o_values_reg[46][13]  (.Q (\o_values[46] [13] ), .CK (n_0_121), .D (sps__n1));
DFF_X1 \o_values_reg[46][14]  (.Q (\o_values[46] [14] ), .CK (n_0_121), .D (sps__n13));
DFF_X1 \o_values_reg[46][15]  (.Q (\o_values[46] [15] ), .CK (n_0_121), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[46]_reg  (.GCK (n_0_121), .CK (clk), .E (n_0_37), .SE (1'b0 ));
DFF_X1 \o_values_reg[47][0]  (.Q (\o_values[47] [0] ), .CK (n_0_120), .D (sps__n16));
DFF_X1 \o_values_reg[47][1]  (.Q (\o_values[47] [1] ), .CK (n_0_120), .D (sps__n25));
DFF_X1 \o_values_reg[47][2]  (.Q (\o_values[47] [2] ), .CK (n_0_120), .D (sps__n19));
DFF_X1 \o_values_reg[47][3]  (.Q (\o_values[47] [3] ), .CK (n_0_120), .D (sps__n28));
DFF_X1 \o_values_reg[47][4]  (.Q (\o_values[47] [4] ), .CK (n_0_120), .D (sps__n31));
DFF_X1 \o_values_reg[47][5]  (.Q (\o_values[47] [5] ), .CK (n_0_120), .D (sps__n34));
DFF_X1 \o_values_reg[47][6]  (.Q (\o_values[47] [6] ), .CK (n_0_120), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[47][7]  (.Q (\o_values[47] [7] ), .CK (n_0_120), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[47][8]  (.Q (\o_values[47] [8] ), .CK (n_0_120), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[47][9]  (.Q (\o_values[47] [9] ), .CK (n_0_120), .D (sps__n37));
DFF_X1 \o_values_reg[47][10]  (.Q (\o_values[47] [10] ), .CK (n_0_120), .D (sps__n4));
DFF_X1 \o_values_reg[47][11]  (.Q (\o_values[47] [11] ), .CK (n_0_120), .D (sps__n10));
DFF_X1 \o_values_reg[47][12]  (.Q (\o_values[47] [12] ), .CK (n_0_120), .D (sps__n7));
DFF_X1 \o_values_reg[47][13]  (.Q (\o_values[47] [13] ), .CK (n_0_120), .D (sps__n1));
DFF_X1 \o_values_reg[47][14]  (.Q (\o_values[47] [14] ), .CK (n_0_120), .D (sps__n13));
DFF_X1 \o_values_reg[47][15]  (.Q (\o_values[47] [15] ), .CK (n_0_120), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[47]_reg  (.GCK (n_0_120), .CK (clk), .E (n_0_36), .SE (1'b0 ));
DFF_X1 \o_values_reg[48][0]  (.Q (\o_values[48] [0] ), .CK (n_0_119), .D (sps__n16));
DFF_X1 \o_values_reg[48][1]  (.Q (\o_values[48] [1] ), .CK (n_0_119), .D (sps__n25));
DFF_X1 \o_values_reg[48][2]  (.Q (\o_values[48] [2] ), .CK (n_0_119), .D (sps__n19));
DFF_X1 \o_values_reg[48][3]  (.Q (\o_values[48] [3] ), .CK (n_0_119), .D (sps__n28));
DFF_X1 \o_values_reg[48][4]  (.Q (\o_values[48] [4] ), .CK (n_0_119), .D (sps__n31));
DFF_X1 \o_values_reg[48][5]  (.Q (\o_values[48] [5] ), .CK (n_0_119), .D (sps__n34));
DFF_X1 \o_values_reg[48][6]  (.Q (\o_values[48] [6] ), .CK (n_0_119), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[48][7]  (.Q (\o_values[48] [7] ), .CK (n_0_119), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[48][8]  (.Q (\o_values[48] [8] ), .CK (n_0_119), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[48][9]  (.Q (\o_values[48] [9] ), .CK (n_0_119), .D (sps__n37));
DFF_X1 \o_values_reg[48][10]  (.Q (\o_values[48] [10] ), .CK (n_0_119), .D (sps__n4));
DFF_X1 \o_values_reg[48][11]  (.Q (\o_values[48] [11] ), .CK (n_0_119), .D (sps__n10));
DFF_X1 \o_values_reg[48][12]  (.Q (\o_values[48] [12] ), .CK (n_0_119), .D (sps__n7));
DFF_X1 \o_values_reg[48][13]  (.Q (\o_values[48] [13] ), .CK (n_0_119), .D (sps__n1));
DFF_X1 \o_values_reg[48][14]  (.Q (\o_values[48] [14] ), .CK (n_0_119), .D (sps__n13));
DFF_X1 \o_values_reg[48][15]  (.Q (\o_values[48] [15] ), .CK (n_0_119), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[48]_reg  (.GCK (n_0_119), .CK (clk), .E (n_0_35), .SE (1'b0 ));
DFF_X1 \o_values_reg[49][0]  (.Q (\o_values[49] [0] ), .CK (n_0_118), .D (sps__n16));
DFF_X1 \o_values_reg[49][1]  (.Q (\o_values[49] [1] ), .CK (n_0_118), .D (sps__n25));
DFF_X1 \o_values_reg[49][2]  (.Q (\o_values[49] [2] ), .CK (n_0_118), .D (sps__n19));
DFF_X1 \o_values_reg[49][3]  (.Q (\o_values[49] [3] ), .CK (n_0_118), .D (sps__n28));
DFF_X1 \o_values_reg[49][4]  (.Q (\o_values[49] [4] ), .CK (n_0_118), .D (sps__n31));
DFF_X1 \o_values_reg[49][5]  (.Q (\o_values[49] [5] ), .CK (n_0_118), .D (sps__n34));
DFF_X1 \o_values_reg[49][6]  (.Q (\o_values[49] [6] ), .CK (n_0_118), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[49][7]  (.Q (\o_values[49] [7] ), .CK (n_0_118), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[49][8]  (.Q (\o_values[49] [8] ), .CK (n_0_118), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[49][9]  (.Q (\o_values[49] [9] ), .CK (n_0_118), .D (sps__n37));
DFF_X1 \o_values_reg[49][10]  (.Q (\o_values[49] [10] ), .CK (n_0_118), .D (sps__n4));
DFF_X1 \o_values_reg[49][11]  (.Q (\o_values[49] [11] ), .CK (n_0_118), .D (sps__n10));
DFF_X1 \o_values_reg[49][12]  (.Q (\o_values[49] [12] ), .CK (n_0_118), .D (sps__n7));
DFF_X1 \o_values_reg[49][13]  (.Q (\o_values[49] [13] ), .CK (n_0_118), .D (sps__n1));
DFF_X1 \o_values_reg[49][14]  (.Q (\o_values[49] [14] ), .CK (n_0_118), .D (sps__n13));
DFF_X1 \o_values_reg[49][15]  (.Q (\o_values[49] [15] ), .CK (n_0_118), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[49]_reg  (.GCK (n_0_118), .CK (clk), .E (n_0_34), .SE (1'b0 ));
DFF_X1 \o_values_reg[50][0]  (.Q (\o_values[50] [0] ), .CK (n_0_117), .D (sps__n16));
DFF_X1 \o_values_reg[50][1]  (.Q (\o_values[50] [1] ), .CK (n_0_117), .D (sps__n25));
DFF_X1 \o_values_reg[50][2]  (.Q (\o_values[50] [2] ), .CK (n_0_117), .D (sps__n19));
DFF_X1 \o_values_reg[50][3]  (.Q (\o_values[50] [3] ), .CK (n_0_117), .D (sps__n28));
DFF_X1 \o_values_reg[50][4]  (.Q (\o_values[50] [4] ), .CK (n_0_117), .D (sps__n31));
DFF_X1 \o_values_reg[50][5]  (.Q (\o_values[50] [5] ), .CK (n_0_117), .D (sps__n34));
DFF_X1 \o_values_reg[50][6]  (.Q (\o_values[50] [6] ), .CK (n_0_117), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[50][7]  (.Q (\o_values[50] [7] ), .CK (n_0_117), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[50][8]  (.Q (\o_values[50] [8] ), .CK (n_0_117), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[50][9]  (.Q (\o_values[50] [9] ), .CK (n_0_117), .D (sps__n37));
DFF_X1 \o_values_reg[50][10]  (.Q (\o_values[50] [10] ), .CK (n_0_117), .D (sps__n4));
DFF_X1 \o_values_reg[50][11]  (.Q (\o_values[50] [11] ), .CK (n_0_117), .D (sps__n10));
DFF_X1 \o_values_reg[50][12]  (.Q (\o_values[50] [12] ), .CK (n_0_117), .D (sps__n7));
DFF_X1 \o_values_reg[50][13]  (.Q (\o_values[50] [13] ), .CK (n_0_117), .D (sps__n1));
DFF_X1 \o_values_reg[50][14]  (.Q (\o_values[50] [14] ), .CK (n_0_117), .D (sps__n13));
DFF_X1 \o_values_reg[50][15]  (.Q (\o_values[50] [15] ), .CK (n_0_117), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[50]_reg  (.GCK (n_0_117), .CK (clk), .E (n_0_33), .SE (1'b0 ));
DFF_X1 \o_values_reg[51][0]  (.Q (\o_values[51] [0] ), .CK (n_0_116), .D (sps__n16));
DFF_X1 \o_values_reg[51][1]  (.Q (\o_values[51] [1] ), .CK (n_0_116), .D (sps__n25));
DFF_X1 \o_values_reg[51][2]  (.Q (\o_values[51] [2] ), .CK (n_0_116), .D (sps__n19));
DFF_X1 \o_values_reg[51][3]  (.Q (\o_values[51] [3] ), .CK (n_0_116), .D (sps__n28));
DFF_X1 \o_values_reg[51][4]  (.Q (\o_values[51] [4] ), .CK (n_0_116), .D (sps__n31));
DFF_X1 \o_values_reg[51][5]  (.Q (\o_values[51] [5] ), .CK (n_0_116), .D (sps__n34));
DFF_X1 \o_values_reg[51][6]  (.Q (\o_values[51] [6] ), .CK (n_0_116), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[51][7]  (.Q (\o_values[51] [7] ), .CK (n_0_116), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[51][8]  (.Q (\o_values[51] [8] ), .CK (n_0_116), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[51][9]  (.Q (\o_values[51] [9] ), .CK (n_0_116), .D (sps__n37));
DFF_X1 \o_values_reg[51][10]  (.Q (\o_values[51] [10] ), .CK (n_0_116), .D (sps__n4));
DFF_X1 \o_values_reg[51][11]  (.Q (\o_values[51] [11] ), .CK (n_0_116), .D (sps__n10));
DFF_X1 \o_values_reg[51][12]  (.Q (\o_values[51] [12] ), .CK (n_0_116), .D (sps__n7));
DFF_X1 \o_values_reg[51][13]  (.Q (\o_values[51] [13] ), .CK (n_0_116), .D (sps__n1));
DFF_X1 \o_values_reg[51][14]  (.Q (\o_values[51] [14] ), .CK (n_0_116), .D (sps__n13));
DFF_X1 \o_values_reg[51][15]  (.Q (\o_values[51] [15] ), .CK (n_0_116), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[51]_reg  (.GCK (n_0_116), .CK (clk), .E (n_0_32), .SE (1'b0 ));
DFF_X1 \o_values_reg[52][0]  (.Q (\o_values[52] [0] ), .CK (n_0_115), .D (sps__n16));
DFF_X1 \o_values_reg[52][1]  (.Q (\o_values[52] [1] ), .CK (n_0_115), .D (sps__n25));
DFF_X1 \o_values_reg[52][2]  (.Q (\o_values[52] [2] ), .CK (n_0_115), .D (sps__n19));
DFF_X1 \o_values_reg[52][3]  (.Q (\o_values[52] [3] ), .CK (n_0_115), .D (sps__n28));
DFF_X1 \o_values_reg[52][4]  (.Q (\o_values[52] [4] ), .CK (n_0_115), .D (sps__n31));
DFF_X1 \o_values_reg[52][5]  (.Q (\o_values[52] [5] ), .CK (n_0_115), .D (sps__n34));
DFF_X1 \o_values_reg[52][6]  (.Q (\o_values[52] [6] ), .CK (n_0_115), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[52][7]  (.Q (\o_values[52] [7] ), .CK (n_0_115), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[52][8]  (.Q (\o_values[52] [8] ), .CK (n_0_115), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[52][9]  (.Q (\o_values[52] [9] ), .CK (n_0_115), .D (sps__n37));
DFF_X1 \o_values_reg[52][10]  (.Q (\o_values[52] [10] ), .CK (n_0_115), .D (sps__n4));
DFF_X1 \o_values_reg[52][11]  (.Q (\o_values[52] [11] ), .CK (n_0_115), .D (sps__n10));
DFF_X1 \o_values_reg[52][12]  (.Q (\o_values[52] [12] ), .CK (n_0_115), .D (sps__n7));
DFF_X1 \o_values_reg[52][13]  (.Q (\o_values[52] [13] ), .CK (n_0_115), .D (sps__n1));
DFF_X1 \o_values_reg[52][14]  (.Q (\o_values[52] [14] ), .CK (n_0_115), .D (sps__n13));
DFF_X1 \o_values_reg[52][15]  (.Q (\o_values[52] [15] ), .CK (n_0_115), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[52]_reg  (.GCK (n_0_115), .CK (clk), .E (n_0_31), .SE (1'b0 ));
DFF_X1 \o_values_reg[53][0]  (.Q (\o_values[53] [0] ), .CK (n_0_114), .D (sps__n16));
DFF_X1 \o_values_reg[53][1]  (.Q (\o_values[53] [1] ), .CK (n_0_114), .D (sps__n25));
DFF_X1 \o_values_reg[53][2]  (.Q (\o_values[53] [2] ), .CK (n_0_114), .D (sps__n19));
DFF_X1 \o_values_reg[53][3]  (.Q (\o_values[53] [3] ), .CK (n_0_114), .D (sps__n28));
DFF_X1 \o_values_reg[53][4]  (.Q (\o_values[53] [4] ), .CK (n_0_114), .D (sps__n31));
DFF_X1 \o_values_reg[53][5]  (.Q (\o_values[53] [5] ), .CK (n_0_114), .D (sps__n34));
DFF_X1 \o_values_reg[53][6]  (.Q (\o_values[53] [6] ), .CK (n_0_114), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[53][7]  (.Q (\o_values[53] [7] ), .CK (n_0_114), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[53][8]  (.Q (\o_values[53] [8] ), .CK (n_0_114), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[53][9]  (.Q (\o_values[53] [9] ), .CK (n_0_114), .D (sps__n37));
DFF_X1 \o_values_reg[53][10]  (.Q (\o_values[53] [10] ), .CK (n_0_114), .D (sps__n4));
DFF_X1 \o_values_reg[53][11]  (.Q (\o_values[53] [11] ), .CK (n_0_114), .D (sps__n10));
DFF_X1 \o_values_reg[53][12]  (.Q (\o_values[53] [12] ), .CK (n_0_114), .D (sps__n7));
DFF_X1 \o_values_reg[53][13]  (.Q (\o_values[53] [13] ), .CK (n_0_114), .D (sps__n1));
DFF_X1 \o_values_reg[53][14]  (.Q (\o_values[53] [14] ), .CK (n_0_114), .D (sps__n13));
DFF_X1 \o_values_reg[53][15]  (.Q (\o_values[53] [15] ), .CK (n_0_114), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[53]_reg  (.GCK (n_0_114), .CK (clk), .E (n_0_30), .SE (1'b0 ));
DFF_X1 \o_values_reg[54][0]  (.Q (\o_values[54] [0] ), .CK (n_0_113), .D (sps__n16));
DFF_X1 \o_values_reg[54][1]  (.Q (\o_values[54] [1] ), .CK (n_0_113), .D (sps__n25));
DFF_X1 \o_values_reg[54][2]  (.Q (\o_values[54] [2] ), .CK (n_0_113), .D (sps__n19));
DFF_X1 \o_values_reg[54][3]  (.Q (\o_values[54] [3] ), .CK (n_0_113), .D (sps__n28));
DFF_X1 \o_values_reg[54][4]  (.Q (\o_values[54] [4] ), .CK (n_0_113), .D (sps__n31));
DFF_X1 \o_values_reg[54][5]  (.Q (\o_values[54] [5] ), .CK (n_0_113), .D (sps__n34));
DFF_X1 \o_values_reg[54][6]  (.Q (\o_values[54] [6] ), .CK (n_0_113), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[54][7]  (.Q (\o_values[54] [7] ), .CK (n_0_113), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[54][8]  (.Q (\o_values[54] [8] ), .CK (n_0_113), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[54][9]  (.Q (\o_values[54] [9] ), .CK (n_0_113), .D (sps__n37));
DFF_X1 \o_values_reg[54][10]  (.Q (\o_values[54] [10] ), .CK (n_0_113), .D (sps__n4));
DFF_X1 \o_values_reg[54][11]  (.Q (\o_values[54] [11] ), .CK (n_0_113), .D (sps__n10));
DFF_X1 \o_values_reg[54][12]  (.Q (\o_values[54] [12] ), .CK (n_0_113), .D (sps__n7));
DFF_X1 \o_values_reg[54][13]  (.Q (\o_values[54] [13] ), .CK (n_0_113), .D (sps__n1));
DFF_X1 \o_values_reg[54][14]  (.Q (\o_values[54] [14] ), .CK (n_0_113), .D (sps__n13));
DFF_X1 \o_values_reg[54][15]  (.Q (\o_values[54] [15] ), .CK (n_0_113), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[54]_reg  (.GCK (n_0_113), .CK (clk), .E (n_0_29), .SE (1'b0 ));
DFF_X1 \o_values_reg[55][0]  (.Q (\o_values[55] [0] ), .CK (n_0_112), .D (sps__n16));
DFF_X1 \o_values_reg[55][1]  (.Q (\o_values[55] [1] ), .CK (n_0_112), .D (sps__n25));
DFF_X1 \o_values_reg[55][2]  (.Q (\o_values[55] [2] ), .CK (n_0_112), .D (sps__n19));
DFF_X1 \o_values_reg[55][3]  (.Q (\o_values[55] [3] ), .CK (n_0_112), .D (sps__n28));
DFF_X1 \o_values_reg[55][4]  (.Q (\o_values[55] [4] ), .CK (n_0_112), .D (sps__n31));
DFF_X1 \o_values_reg[55][5]  (.Q (\o_values[55] [5] ), .CK (n_0_112), .D (sps__n34));
DFF_X1 \o_values_reg[55][6]  (.Q (\o_values[55] [6] ), .CK (n_0_112), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[55][7]  (.Q (\o_values[55] [7] ), .CK (n_0_112), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[55][8]  (.Q (\o_values[55] [8] ), .CK (n_0_112), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[55][9]  (.Q (\o_values[55] [9] ), .CK (n_0_112), .D (sps__n37));
DFF_X1 \o_values_reg[55][10]  (.Q (\o_values[55] [10] ), .CK (n_0_112), .D (sps__n4));
DFF_X1 \o_values_reg[55][11]  (.Q (\o_values[55] [11] ), .CK (n_0_112), .D (sps__n10));
DFF_X1 \o_values_reg[55][12]  (.Q (\o_values[55] [12] ), .CK (n_0_112), .D (sps__n7));
DFF_X1 \o_values_reg[55][13]  (.Q (\o_values[55] [13] ), .CK (n_0_112), .D (sps__n1));
DFF_X1 \o_values_reg[55][14]  (.Q (\o_values[55] [14] ), .CK (n_0_112), .D (sps__n13));
DFF_X1 \o_values_reg[55][15]  (.Q (\o_values[55] [15] ), .CK (n_0_112), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[55]_reg  (.GCK (n_0_112), .CK (clk), .E (n_0_28), .SE (1'b0 ));
DFF_X1 \o_values_reg[56][0]  (.Q (\o_values[56] [0] ), .CK (n_0_111), .D (sps__n16));
DFF_X1 \o_values_reg[56][1]  (.Q (\o_values[56] [1] ), .CK (n_0_111), .D (sps__n25));
DFF_X1 \o_values_reg[56][2]  (.Q (\o_values[56] [2] ), .CK (n_0_111), .D (sps__n19));
DFF_X1 \o_values_reg[56][3]  (.Q (\o_values[56] [3] ), .CK (n_0_111), .D (sps__n28));
DFF_X1 \o_values_reg[56][4]  (.Q (\o_values[56] [4] ), .CK (n_0_111), .D (sps__n31));
DFF_X1 \o_values_reg[56][5]  (.Q (\o_values[56] [5] ), .CK (n_0_111), .D (sps__n34));
DFF_X1 \o_values_reg[56][6]  (.Q (\o_values[56] [6] ), .CK (n_0_111), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[56][7]  (.Q (\o_values[56] [7] ), .CK (n_0_111), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[56][8]  (.Q (\o_values[56] [8] ), .CK (n_0_111), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[56][9]  (.Q (\o_values[56] [9] ), .CK (n_0_111), .D (sps__n37));
DFF_X1 \o_values_reg[56][10]  (.Q (\o_values[56] [10] ), .CK (n_0_111), .D (sps__n4));
DFF_X1 \o_values_reg[56][11]  (.Q (\o_values[56] [11] ), .CK (n_0_111), .D (sps__n10));
DFF_X1 \o_values_reg[56][12]  (.Q (\o_values[56] [12] ), .CK (n_0_111), .D (sps__n7));
DFF_X1 \o_values_reg[56][13]  (.Q (\o_values[56] [13] ), .CK (n_0_111), .D (sps__n1));
DFF_X1 \o_values_reg[56][14]  (.Q (\o_values[56] [14] ), .CK (n_0_111), .D (sps__n13));
DFF_X1 \o_values_reg[56][15]  (.Q (\o_values[56] [15] ), .CK (n_0_111), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[56]_reg  (.GCK (n_0_111), .CK (clk), .E (n_0_27), .SE (1'b0 ));
DFF_X1 \o_values_reg[57][0]  (.Q (\o_values[57] [0] ), .CK (n_0_110), .D (sps__n16));
DFF_X1 \o_values_reg[57][1]  (.Q (\o_values[57] [1] ), .CK (n_0_110), .D (sps__n25));
DFF_X1 \o_values_reg[57][2]  (.Q (\o_values[57] [2] ), .CK (n_0_110), .D (sps__n19));
DFF_X1 \o_values_reg[57][3]  (.Q (\o_values[57] [3] ), .CK (n_0_110), .D (sps__n28));
DFF_X1 \o_values_reg[57][4]  (.Q (\o_values[57] [4] ), .CK (n_0_110), .D (sps__n31));
DFF_X1 \o_values_reg[57][5]  (.Q (\o_values[57] [5] ), .CK (n_0_110), .D (sps__n34));
DFF_X1 \o_values_reg[57][6]  (.Q (\o_values[57] [6] ), .CK (n_0_110), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[57][7]  (.Q (\o_values[57] [7] ), .CK (n_0_110), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[57][8]  (.Q (\o_values[57] [8] ), .CK (n_0_110), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[57][9]  (.Q (\o_values[57] [9] ), .CK (n_0_110), .D (sps__n37));
DFF_X1 \o_values_reg[57][10]  (.Q (\o_values[57] [10] ), .CK (n_0_110), .D (sps__n4));
DFF_X1 \o_values_reg[57][11]  (.Q (\o_values[57] [11] ), .CK (n_0_110), .D (sps__n10));
DFF_X1 \o_values_reg[57][12]  (.Q (\o_values[57] [12] ), .CK (n_0_110), .D (sps__n7));
DFF_X1 \o_values_reg[57][13]  (.Q (\o_values[57] [13] ), .CK (n_0_110), .D (sps__n1));
DFF_X1 \o_values_reg[57][14]  (.Q (\o_values[57] [14] ), .CK (n_0_110), .D (sps__n13));
DFF_X1 \o_values_reg[57][15]  (.Q (\o_values[57] [15] ), .CK (n_0_110), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[57]_reg  (.GCK (n_0_110), .CK (clk), .E (n_0_26), .SE (1'b0 ));
DFF_X1 \o_values_reg[58][0]  (.Q (\o_values[58] [0] ), .CK (n_0_109), .D (sps__n16));
DFF_X1 \o_values_reg[58][1]  (.Q (\o_values[58] [1] ), .CK (n_0_109), .D (sps__n25));
DFF_X1 \o_values_reg[58][2]  (.Q (\o_values[58] [2] ), .CK (n_0_109), .D (sps__n19));
DFF_X1 \o_values_reg[58][3]  (.Q (\o_values[58] [3] ), .CK (n_0_109), .D (sps__n28));
DFF_X1 \o_values_reg[58][4]  (.Q (\o_values[58] [4] ), .CK (n_0_109), .D (sps__n31));
DFF_X1 \o_values_reg[58][5]  (.Q (\o_values[58] [5] ), .CK (n_0_109), .D (sps__n34));
DFF_X1 \o_values_reg[58][6]  (.Q (\o_values[58] [6] ), .CK (n_0_109), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[58][7]  (.Q (\o_values[58] [7] ), .CK (n_0_109), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[58][8]  (.Q (\o_values[58] [8] ), .CK (n_0_109), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[58][9]  (.Q (\o_values[58] [9] ), .CK (n_0_109), .D (sps__n37));
DFF_X1 \o_values_reg[58][10]  (.Q (\o_values[58] [10] ), .CK (n_0_109), .D (sps__n4));
DFF_X1 \o_values_reg[58][11]  (.Q (\o_values[58] [11] ), .CK (n_0_109), .D (sps__n10));
DFF_X1 \o_values_reg[58][12]  (.Q (\o_values[58] [12] ), .CK (n_0_109), .D (sps__n7));
DFF_X1 \o_values_reg[58][13]  (.Q (\o_values[58] [13] ), .CK (n_0_109), .D (sps__n1));
DFF_X1 \o_values_reg[58][14]  (.Q (\o_values[58] [14] ), .CK (n_0_109), .D (sps__n13));
DFF_X1 \o_values_reg[58][15]  (.Q (\o_values[58] [15] ), .CK (n_0_109), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[58]_reg  (.GCK (n_0_109), .CK (clk), .E (n_0_25), .SE (1'b0 ));
DFF_X1 \o_values_reg[59][0]  (.Q (\o_values[59] [0] ), .CK (n_0_108), .D (sps__n16));
DFF_X1 \o_values_reg[59][1]  (.Q (\o_values[59] [1] ), .CK (n_0_108), .D (sps__n25));
DFF_X1 \o_values_reg[59][2]  (.Q (\o_values[59] [2] ), .CK (n_0_108), .D (sps__n19));
DFF_X1 \o_values_reg[59][3]  (.Q (\o_values[59] [3] ), .CK (n_0_108), .D (sps__n28));
DFF_X1 \o_values_reg[59][4]  (.Q (\o_values[59] [4] ), .CK (n_0_108), .D (sps__n31));
DFF_X1 \o_values_reg[59][5]  (.Q (\o_values[59] [5] ), .CK (n_0_108), .D (sps__n34));
DFF_X1 \o_values_reg[59][6]  (.Q (\o_values[59] [6] ), .CK (n_0_108), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[59][7]  (.Q (\o_values[59] [7] ), .CK (n_0_108), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[59][8]  (.Q (\o_values[59] [8] ), .CK (n_0_108), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[59][9]  (.Q (\o_values[59] [9] ), .CK (n_0_108), .D (sps__n37));
DFF_X1 \o_values_reg[59][10]  (.Q (\o_values[59] [10] ), .CK (n_0_108), .D (sps__n4));
DFF_X1 \o_values_reg[59][11]  (.Q (\o_values[59] [11] ), .CK (n_0_108), .D (sps__n10));
DFF_X1 \o_values_reg[59][12]  (.Q (\o_values[59] [12] ), .CK (n_0_108), .D (sps__n7));
DFF_X1 \o_values_reg[59][13]  (.Q (\o_values[59] [13] ), .CK (n_0_108), .D (sps__n1));
DFF_X1 \o_values_reg[59][14]  (.Q (\o_values[59] [14] ), .CK (n_0_108), .D (sps__n13));
DFF_X1 \o_values_reg[59][15]  (.Q (\o_values[59] [15] ), .CK (n_0_108), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[59]_reg  (.GCK (n_0_108), .CK (clk), .E (n_0_24), .SE (1'b0 ));
DFF_X1 \o_values_reg[60][0]  (.Q (\o_values[60] [0] ), .CK (n_0_107), .D (sps__n16));
DFF_X1 \o_values_reg[60][1]  (.Q (\o_values[60] [1] ), .CK (n_0_107), .D (sps__n25));
DFF_X1 \o_values_reg[60][2]  (.Q (\o_values[60] [2] ), .CK (n_0_107), .D (sps__n19));
DFF_X1 \o_values_reg[60][3]  (.Q (\o_values[60] [3] ), .CK (n_0_107), .D (sps__n28));
DFF_X1 \o_values_reg[60][4]  (.Q (\o_values[60] [4] ), .CK (n_0_107), .D (sps__n31));
DFF_X1 \o_values_reg[60][5]  (.Q (\o_values[60] [5] ), .CK (n_0_107), .D (sps__n34));
DFF_X1 \o_values_reg[60][6]  (.Q (\o_values[60] [6] ), .CK (n_0_107), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[60][7]  (.Q (\o_values[60] [7] ), .CK (n_0_107), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[60][8]  (.Q (\o_values[60] [8] ), .CK (n_0_107), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[60][9]  (.Q (\o_values[60] [9] ), .CK (n_0_107), .D (sps__n37));
DFF_X1 \o_values_reg[60][10]  (.Q (\o_values[60] [10] ), .CK (n_0_107), .D (sps__n4));
DFF_X1 \o_values_reg[60][11]  (.Q (\o_values[60] [11] ), .CK (n_0_107), .D (sps__n10));
DFF_X1 \o_values_reg[60][12]  (.Q (\o_values[60] [12] ), .CK (n_0_107), .D (sps__n7));
DFF_X1 \o_values_reg[60][13]  (.Q (\o_values[60] [13] ), .CK (n_0_107), .D (sps__n1));
DFF_X1 \o_values_reg[60][14]  (.Q (\o_values[60] [14] ), .CK (n_0_107), .D (sps__n13));
DFF_X1 \o_values_reg[60][15]  (.Q (\o_values[60] [15] ), .CK (n_0_107), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[60]_reg  (.GCK (n_0_107), .CK (clk), .E (n_0_23), .SE (1'b0 ));
DFF_X1 \o_values_reg[61][0]  (.Q (\o_values[61] [0] ), .CK (n_0_106), .D (sps__n16));
DFF_X1 \o_values_reg[61][1]  (.Q (\o_values[61] [1] ), .CK (n_0_106), .D (sps__n25));
DFF_X1 \o_values_reg[61][2]  (.Q (\o_values[61] [2] ), .CK (n_0_106), .D (sps__n19));
DFF_X1 \o_values_reg[61][3]  (.Q (\o_values[61] [3] ), .CK (n_0_106), .D (sps__n28));
DFF_X1 \o_values_reg[61][4]  (.Q (\o_values[61] [4] ), .CK (n_0_106), .D (sps__n31));
DFF_X1 \o_values_reg[61][5]  (.Q (\o_values[61] [5] ), .CK (n_0_106), .D (sps__n34));
DFF_X1 \o_values_reg[61][6]  (.Q (\o_values[61] [6] ), .CK (n_0_106), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[61][7]  (.Q (\o_values[61] [7] ), .CK (n_0_106), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[61][8]  (.Q (\o_values[61] [8] ), .CK (n_0_106), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[61][9]  (.Q (\o_values[61] [9] ), .CK (n_0_106), .D (sps__n37));
DFF_X1 \o_values_reg[61][10]  (.Q (\o_values[61] [10] ), .CK (n_0_106), .D (sps__n4));
DFF_X1 \o_values_reg[61][11]  (.Q (\o_values[61] [11] ), .CK (n_0_106), .D (sps__n10));
DFF_X1 \o_values_reg[61][12]  (.Q (\o_values[61] [12] ), .CK (n_0_106), .D (sps__n7));
DFF_X1 \o_values_reg[61][13]  (.Q (\o_values[61] [13] ), .CK (n_0_106), .D (sps__n1));
DFF_X1 \o_values_reg[61][14]  (.Q (\o_values[61] [14] ), .CK (n_0_106), .D (sps__n13));
DFF_X1 \o_values_reg[61][15]  (.Q (\o_values[61] [15] ), .CK (n_0_106), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[61]_reg  (.GCK (n_0_106), .CK (clk), .E (n_0_22), .SE (1'b0 ));
DFF_X1 \o_values_reg[62][0]  (.Q (\o_values[62] [0] ), .CK (n_0_105), .D (sps__n16));
DFF_X1 \o_values_reg[62][1]  (.Q (\o_values[62] [1] ), .CK (n_0_105), .D (sps__n25));
DFF_X1 \o_values_reg[62][2]  (.Q (\o_values[62] [2] ), .CK (n_0_105), .D (sps__n19));
DFF_X1 \o_values_reg[62][3]  (.Q (\o_values[62] [3] ), .CK (n_0_105), .D (sps__n28));
DFF_X1 \o_values_reg[62][4]  (.Q (\o_values[62] [4] ), .CK (n_0_105), .D (sps__n31));
DFF_X1 \o_values_reg[62][5]  (.Q (\o_values[62] [5] ), .CK (n_0_105), .D (sps__n34));
DFF_X1 \o_values_reg[62][6]  (.Q (\o_values[62] [6] ), .CK (n_0_105), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[62][7]  (.Q (\o_values[62] [7] ), .CK (n_0_105), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[62][8]  (.Q (\o_values[62] [8] ), .CK (n_0_105), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[62][9]  (.Q (\o_values[62] [9] ), .CK (n_0_105), .D (sps__n37));
DFF_X1 \o_values_reg[62][10]  (.Q (\o_values[62] [10] ), .CK (n_0_105), .D (sps__n4));
DFF_X1 \o_values_reg[62][11]  (.Q (\o_values[62] [11] ), .CK (n_0_105), .D (sps__n10));
DFF_X1 \o_values_reg[62][12]  (.Q (\o_values[62] [12] ), .CK (n_0_105), .D (sps__n7));
DFF_X1 \o_values_reg[62][13]  (.Q (\o_values[62] [13] ), .CK (n_0_105), .D (sps__n1));
DFF_X1 \o_values_reg[62][14]  (.Q (\o_values[62] [14] ), .CK (n_0_105), .D (sps__n13));
DFF_X1 \o_values_reg[62][15]  (.Q (\o_values[62] [15] ), .CK (n_0_105), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[62]_reg  (.GCK (n_0_105), .CK (clk), .E (n_0_21), .SE (1'b0 ));
DFF_X1 \o_values_reg[63][0]  (.Q (\o_values[63] [0] ), .CK (n_0_104), .D (sps__n16));
DFF_X1 \o_values_reg[63][1]  (.Q (\o_values[63] [1] ), .CK (n_0_104), .D (sps__n25));
DFF_X1 \o_values_reg[63][2]  (.Q (\o_values[63] [2] ), .CK (n_0_104), .D (sps__n19));
DFF_X1 \o_values_reg[63][3]  (.Q (\o_values[63] [3] ), .CK (n_0_104), .D (sps__n28));
DFF_X1 \o_values_reg[63][4]  (.Q (\o_values[63] [4] ), .CK (n_0_104), .D (sps__n31));
DFF_X1 \o_values_reg[63][5]  (.Q (\o_values[63] [5] ), .CK (n_0_104), .D (sps__n34));
DFF_X1 \o_values_reg[63][6]  (.Q (\o_values[63] [6] ), .CK (n_0_104), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[63][7]  (.Q (\o_values[63] [7] ), .CK (n_0_104), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[63][8]  (.Q (\o_values[63] [8] ), .CK (n_0_104), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[63][9]  (.Q (\o_values[63] [9] ), .CK (n_0_104), .D (sps__n37));
DFF_X1 \o_values_reg[63][10]  (.Q (\o_values[63] [10] ), .CK (n_0_104), .D (sps__n4));
DFF_X1 \o_values_reg[63][11]  (.Q (\o_values[63] [11] ), .CK (n_0_104), .D (sps__n10));
DFF_X1 \o_values_reg[63][12]  (.Q (\o_values[63] [12] ), .CK (n_0_104), .D (sps__n7));
DFF_X1 \o_values_reg[63][13]  (.Q (\o_values[63] [13] ), .CK (n_0_104), .D (sps__n1));
DFF_X1 \o_values_reg[63][14]  (.Q (\o_values[63] [14] ), .CK (n_0_104), .D (sps__n13));
DFF_X1 \o_values_reg[63][15]  (.Q (\o_values[63] [15] ), .CK (n_0_104), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[63]_reg  (.GCK (n_0_104), .CK (clk), .E (n_0_20), .SE (1'b0 ));
DFF_X1 \o_values_reg[64][0]  (.Q (\o_values[64] [0] ), .CK (n_0_103), .D (sps__n16));
DFF_X1 \o_values_reg[64][1]  (.Q (\o_values[64] [1] ), .CK (n_0_103), .D (sps__n25));
DFF_X1 \o_values_reg[64][2]  (.Q (\o_values[64] [2] ), .CK (n_0_103), .D (sps__n19));
DFF_X1 \o_values_reg[64][3]  (.Q (\o_values[64] [3] ), .CK (n_0_103), .D (sps__n28));
DFF_X1 \o_values_reg[64][4]  (.Q (\o_values[64] [4] ), .CK (n_0_103), .D (sps__n31));
DFF_X1 \o_values_reg[64][5]  (.Q (\o_values[64] [5] ), .CK (n_0_103), .D (sps__n34));
DFF_X1 \o_values_reg[64][6]  (.Q (\o_values[64] [6] ), .CK (n_0_103), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[64][7]  (.Q (\o_values[64] [7] ), .CK (n_0_103), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[64][8]  (.Q (\o_values[64] [8] ), .CK (n_0_103), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[64][9]  (.Q (\o_values[64] [9] ), .CK (n_0_103), .D (sps__n37));
DFF_X1 \o_values_reg[64][10]  (.Q (\o_values[64] [10] ), .CK (n_0_103), .D (sps__n4));
DFF_X1 \o_values_reg[64][11]  (.Q (\o_values[64] [11] ), .CK (n_0_103), .D (sps__n10));
DFF_X1 \o_values_reg[64][12]  (.Q (\o_values[64] [12] ), .CK (n_0_103), .D (sps__n7));
DFF_X1 \o_values_reg[64][13]  (.Q (\o_values[64] [13] ), .CK (n_0_103), .D (sps__n1));
DFF_X1 \o_values_reg[64][14]  (.Q (\o_values[64] [14] ), .CK (n_0_103), .D (sps__n13));
DFF_X1 \o_values_reg[64][15]  (.Q (\o_values[64] [15] ), .CK (n_0_103), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[64]_reg  (.GCK (n_0_103), .CK (clk), .E (n_0_19), .SE (1'b0 ));
DFF_X1 \o_values_reg[65][0]  (.Q (\o_values[65] [0] ), .CK (n_0_102), .D (sps__n16));
DFF_X1 \o_values_reg[65][1]  (.Q (\o_values[65] [1] ), .CK (n_0_102), .D (sps__n25));
DFF_X1 \o_values_reg[65][2]  (.Q (\o_values[65] [2] ), .CK (n_0_102), .D (sps__n19));
DFF_X1 \o_values_reg[65][3]  (.Q (\o_values[65] [3] ), .CK (n_0_102), .D (sps__n28));
DFF_X1 \o_values_reg[65][4]  (.Q (\o_values[65] [4] ), .CK (n_0_102), .D (sps__n31));
DFF_X1 \o_values_reg[65][5]  (.Q (\o_values[65] [5] ), .CK (n_0_102), .D (sps__n34));
DFF_X1 \o_values_reg[65][6]  (.Q (\o_values[65] [6] ), .CK (n_0_102), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[65][7]  (.Q (\o_values[65] [7] ), .CK (n_0_102), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[65][8]  (.Q (\o_values[65] [8] ), .CK (n_0_102), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[65][9]  (.Q (\o_values[65] [9] ), .CK (n_0_102), .D (sps__n37));
DFF_X1 \o_values_reg[65][10]  (.Q (\o_values[65] [10] ), .CK (n_0_102), .D (sps__n4));
DFF_X1 \o_values_reg[65][11]  (.Q (\o_values[65] [11] ), .CK (n_0_102), .D (sps__n10));
DFF_X1 \o_values_reg[65][12]  (.Q (\o_values[65] [12] ), .CK (n_0_102), .D (sps__n7));
DFF_X1 \o_values_reg[65][13]  (.Q (\o_values[65] [13] ), .CK (n_0_102), .D (sps__n1));
DFF_X1 \o_values_reg[65][14]  (.Q (\o_values[65] [14] ), .CK (n_0_102), .D (sps__n13));
DFF_X1 \o_values_reg[65][15]  (.Q (\o_values[65] [15] ), .CK (n_0_102), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[65]_reg  (.GCK (n_0_102), .CK (clk), .E (n_0_18), .SE (1'b0 ));
DFF_X1 \o_values_reg[66][0]  (.Q (\o_values[66] [0] ), .CK (n_0_101), .D (sps__n16));
DFF_X1 \o_values_reg[66][1]  (.Q (\o_values[66] [1] ), .CK (n_0_101), .D (sps__n25));
DFF_X1 \o_values_reg[66][2]  (.Q (\o_values[66] [2] ), .CK (n_0_101), .D (sps__n19));
DFF_X1 \o_values_reg[66][3]  (.Q (\o_values[66] [3] ), .CK (n_0_101), .D (sps__n28));
DFF_X1 \o_values_reg[66][4]  (.Q (\o_values[66] [4] ), .CK (n_0_101), .D (sps__n31));
DFF_X1 \o_values_reg[66][5]  (.Q (\o_values[66] [5] ), .CK (n_0_101), .D (sps__n34));
DFF_X1 \o_values_reg[66][6]  (.Q (\o_values[66] [6] ), .CK (n_0_101), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[66][7]  (.Q (\o_values[66] [7] ), .CK (n_0_101), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[66][8]  (.Q (\o_values[66] [8] ), .CK (n_0_101), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[66][9]  (.Q (\o_values[66] [9] ), .CK (n_0_101), .D (sps__n37));
DFF_X1 \o_values_reg[66][10]  (.Q (\o_values[66] [10] ), .CK (n_0_101), .D (sps__n4));
DFF_X1 \o_values_reg[66][11]  (.Q (\o_values[66] [11] ), .CK (n_0_101), .D (sps__n10));
DFF_X1 \o_values_reg[66][12]  (.Q (\o_values[66] [12] ), .CK (n_0_101), .D (sps__n7));
DFF_X1 \o_values_reg[66][13]  (.Q (\o_values[66] [13] ), .CK (n_0_101), .D (sps__n1));
DFF_X1 \o_values_reg[66][14]  (.Q (\o_values[66] [14] ), .CK (n_0_101), .D (sps__n13));
DFF_X1 \o_values_reg[66][15]  (.Q (\o_values[66] [15] ), .CK (n_0_101), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[66]_reg  (.GCK (n_0_101), .CK (clk), .E (n_0_17), .SE (1'b0 ));
DFF_X1 \o_values_reg[67][0]  (.Q (\o_values[67] [0] ), .CK (n_0_100), .D (sps__n16));
DFF_X1 \o_values_reg[67][1]  (.Q (\o_values[67] [1] ), .CK (n_0_100), .D (sps__n25));
DFF_X1 \o_values_reg[67][2]  (.Q (\o_values[67] [2] ), .CK (n_0_100), .D (sps__n19));
DFF_X1 \o_values_reg[67][3]  (.Q (\o_values[67] [3] ), .CK (n_0_100), .D (sps__n28));
DFF_X1 \o_values_reg[67][4]  (.Q (\o_values[67] [4] ), .CK (n_0_100), .D (sps__n31));
DFF_X1 \o_values_reg[67][5]  (.Q (\o_values[67] [5] ), .CK (n_0_100), .D (sps__n34));
DFF_X1 \o_values_reg[67][6]  (.Q (\o_values[67] [6] ), .CK (n_0_100), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[67][7]  (.Q (\o_values[67] [7] ), .CK (n_0_100), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[67][8]  (.Q (\o_values[67] [8] ), .CK (n_0_100), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[67][9]  (.Q (\o_values[67] [9] ), .CK (n_0_100), .D (sps__n37));
DFF_X1 \o_values_reg[67][10]  (.Q (\o_values[67] [10] ), .CK (n_0_100), .D (sps__n4));
DFF_X1 \o_values_reg[67][11]  (.Q (\o_values[67] [11] ), .CK (n_0_100), .D (sps__n10));
DFF_X1 \o_values_reg[67][12]  (.Q (\o_values[67] [12] ), .CK (n_0_100), .D (sps__n7));
DFF_X1 \o_values_reg[67][13]  (.Q (\o_values[67] [13] ), .CK (n_0_100), .D (sps__n1));
DFF_X1 \o_values_reg[67][14]  (.Q (\o_values[67] [14] ), .CK (n_0_100), .D (sps__n13));
DFF_X1 \o_values_reg[67][15]  (.Q (\o_values[67] [15] ), .CK (n_0_100), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[67]_reg  (.GCK (n_0_100), .CK (clk), .E (n_0_16), .SE (1'b0 ));
DFF_X1 \o_values_reg[68][0]  (.Q (\o_values[68] [0] ), .CK (n_0_99), .D (sps__n16));
DFF_X1 \o_values_reg[68][1]  (.Q (\o_values[68] [1] ), .CK (n_0_99), .D (sps__n25));
DFF_X1 \o_values_reg[68][2]  (.Q (\o_values[68] [2] ), .CK (n_0_99), .D (sps__n19));
DFF_X1 \o_values_reg[68][3]  (.Q (\o_values[68] [3] ), .CK (n_0_99), .D (sps__n28));
DFF_X1 \o_values_reg[68][4]  (.Q (\o_values[68] [4] ), .CK (n_0_99), .D (sps__n31));
DFF_X1 \o_values_reg[68][5]  (.Q (\o_values[68] [5] ), .CK (n_0_99), .D (sps__n34));
DFF_X1 \o_values_reg[68][6]  (.Q (\o_values[68] [6] ), .CK (n_0_99), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[68][7]  (.Q (\o_values[68] [7] ), .CK (n_0_99), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[68][8]  (.Q (\o_values[68] [8] ), .CK (n_0_99), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[68][9]  (.Q (\o_values[68] [9] ), .CK (n_0_99), .D (sps__n37));
DFF_X1 \o_values_reg[68][10]  (.Q (\o_values[68] [10] ), .CK (n_0_99), .D (sps__n4));
DFF_X1 \o_values_reg[68][11]  (.Q (\o_values[68] [11] ), .CK (n_0_99), .D (sps__n10));
DFF_X1 \o_values_reg[68][12]  (.Q (\o_values[68] [12] ), .CK (n_0_99), .D (sps__n7));
DFF_X1 \o_values_reg[68][13]  (.Q (\o_values[68] [13] ), .CK (n_0_99), .D (sps__n1));
DFF_X1 \o_values_reg[68][14]  (.Q (\o_values[68] [14] ), .CK (n_0_99), .D (sps__n13));
DFF_X1 \o_values_reg[68][15]  (.Q (\o_values[68] [15] ), .CK (n_0_99), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[68]_reg  (.GCK (n_0_99), .CK (clk), .E (n_0_15), .SE (1'b0 ));
DFF_X1 \o_values_reg[69][0]  (.Q (\o_values[69] [0] ), .CK (n_0_98), .D (sps__n16));
DFF_X1 \o_values_reg[69][1]  (.Q (\o_values[69] [1] ), .CK (n_0_98), .D (sps__n25));
DFF_X1 \o_values_reg[69][2]  (.Q (\o_values[69] [2] ), .CK (n_0_98), .D (sps__n19));
DFF_X1 \o_values_reg[69][3]  (.Q (\o_values[69] [3] ), .CK (n_0_98), .D (sps__n28));
DFF_X1 \o_values_reg[69][4]  (.Q (\o_values[69] [4] ), .CK (n_0_98), .D (sps__n31));
DFF_X1 \o_values_reg[69][5]  (.Q (\o_values[69] [5] ), .CK (n_0_98), .D (sps__n34));
DFF_X1 \o_values_reg[69][6]  (.Q (\o_values[69] [6] ), .CK (n_0_98), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[69][7]  (.Q (\o_values[69] [7] ), .CK (n_0_98), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[69][8]  (.Q (\o_values[69] [8] ), .CK (n_0_98), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[69][9]  (.Q (\o_values[69] [9] ), .CK (n_0_98), .D (sps__n37));
DFF_X1 \o_values_reg[69][10]  (.Q (\o_values[69] [10] ), .CK (n_0_98), .D (sps__n4));
DFF_X1 \o_values_reg[69][11]  (.Q (\o_values[69] [11] ), .CK (n_0_98), .D (sps__n10));
DFF_X1 \o_values_reg[69][12]  (.Q (\o_values[69] [12] ), .CK (n_0_98), .D (sps__n7));
DFF_X1 \o_values_reg[69][13]  (.Q (\o_values[69] [13] ), .CK (n_0_98), .D (sps__n1));
DFF_X1 \o_values_reg[69][14]  (.Q (\o_values[69] [14] ), .CK (n_0_98), .D (sps__n13));
DFF_X1 \o_values_reg[69][15]  (.Q (\o_values[69] [15] ), .CK (n_0_98), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[69]_reg  (.GCK (n_0_98), .CK (clk), .E (n_0_14), .SE (1'b0 ));
DFF_X1 \o_values_reg[70][0]  (.Q (\o_values[70] [0] ), .CK (n_0_97), .D (sps__n16));
DFF_X1 \o_values_reg[70][1]  (.Q (\o_values[70] [1] ), .CK (n_0_97), .D (sps__n25));
DFF_X1 \o_values_reg[70][2]  (.Q (\o_values[70] [2] ), .CK (n_0_97), .D (sps__n19));
DFF_X1 \o_values_reg[70][3]  (.Q (\o_values[70] [3] ), .CK (n_0_97), .D (sps__n28));
DFF_X1 \o_values_reg[70][4]  (.Q (\o_values[70] [4] ), .CK (n_0_97), .D (sps__n31));
DFF_X1 \o_values_reg[70][5]  (.Q (\o_values[70] [5] ), .CK (n_0_97), .D (sps__n34));
DFF_X1 \o_values_reg[70][6]  (.Q (\o_values[70] [6] ), .CK (n_0_97), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[70][7]  (.Q (\o_values[70] [7] ), .CK (n_0_97), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[70][8]  (.Q (\o_values[70] [8] ), .CK (n_0_97), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[70][9]  (.Q (\o_values[70] [9] ), .CK (n_0_97), .D (sps__n37));
DFF_X1 \o_values_reg[70][10]  (.Q (\o_values[70] [10] ), .CK (n_0_97), .D (sps__n4));
DFF_X1 \o_values_reg[70][11]  (.Q (\o_values[70] [11] ), .CK (n_0_97), .D (sps__n10));
DFF_X1 \o_values_reg[70][12]  (.Q (\o_values[70] [12] ), .CK (n_0_97), .D (sps__n7));
DFF_X1 \o_values_reg[70][13]  (.Q (\o_values[70] [13] ), .CK (n_0_97), .D (sps__n1));
DFF_X1 \o_values_reg[70][14]  (.Q (\o_values[70] [14] ), .CK (n_0_97), .D (sps__n13));
DFF_X1 \o_values_reg[70][15]  (.Q (\o_values[70] [15] ), .CK (n_0_97), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[70]_reg  (.GCK (n_0_97), .CK (clk), .E (n_0_13), .SE (1'b0 ));
DFF_X1 \o_values_reg[71][0]  (.Q (\o_values[71] [0] ), .CK (n_0_96), .D (sps__n16));
DFF_X1 \o_values_reg[71][1]  (.Q (\o_values[71] [1] ), .CK (n_0_96), .D (sps__n25));
DFF_X1 \o_values_reg[71][2]  (.Q (\o_values[71] [2] ), .CK (n_0_96), .D (sps__n19));
DFF_X1 \o_values_reg[71][3]  (.Q (\o_values[71] [3] ), .CK (n_0_96), .D (sps__n28));
DFF_X1 \o_values_reg[71][4]  (.Q (\o_values[71] [4] ), .CK (n_0_96), .D (sps__n31));
DFF_X1 \o_values_reg[71][5]  (.Q (\o_values[71] [5] ), .CK (n_0_96), .D (sps__n34));
DFF_X1 \o_values_reg[71][6]  (.Q (\o_values[71] [6] ), .CK (n_0_96), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[71][7]  (.Q (\o_values[71] [7] ), .CK (n_0_96), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[71][8]  (.Q (\o_values[71] [8] ), .CK (n_0_96), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[71][9]  (.Q (\o_values[71] [9] ), .CK (n_0_96), .D (sps__n37));
DFF_X1 \o_values_reg[71][10]  (.Q (\o_values[71] [10] ), .CK (n_0_96), .D (sps__n4));
DFF_X1 \o_values_reg[71][11]  (.Q (\o_values[71] [11] ), .CK (n_0_96), .D (sps__n10));
DFF_X1 \o_values_reg[71][12]  (.Q (\o_values[71] [12] ), .CK (n_0_96), .D (sps__n7));
DFF_X1 \o_values_reg[71][13]  (.Q (\o_values[71] [13] ), .CK (n_0_96), .D (sps__n1));
DFF_X1 \o_values_reg[71][14]  (.Q (\o_values[71] [14] ), .CK (n_0_96), .D (sps__n13));
DFF_X1 \o_values_reg[71][15]  (.Q (\o_values[71] [15] ), .CK (n_0_96), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[71]_reg  (.GCK (n_0_96), .CK (clk), .E (n_0_12), .SE (1'b0 ));
DFF_X1 \o_values_reg[72][0]  (.Q (\o_values[72] [0] ), .CK (n_0_95), .D (sps__n16));
DFF_X1 \o_values_reg[72][1]  (.Q (\o_values[72] [1] ), .CK (n_0_95), .D (sps__n25));
DFF_X1 \o_values_reg[72][2]  (.Q (\o_values[72] [2] ), .CK (n_0_95), .D (sps__n19));
DFF_X1 \o_values_reg[72][3]  (.Q (\o_values[72] [3] ), .CK (n_0_95), .D (sps__n28));
DFF_X1 \o_values_reg[72][4]  (.Q (\o_values[72] [4] ), .CK (n_0_95), .D (sps__n31));
DFF_X1 \o_values_reg[72][5]  (.Q (\o_values[72] [5] ), .CK (n_0_95), .D (sps__n34));
DFF_X1 \o_values_reg[72][6]  (.Q (\o_values[72] [6] ), .CK (n_0_95), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[72][7]  (.Q (\o_values[72] [7] ), .CK (n_0_95), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[72][8]  (.Q (\o_values[72] [8] ), .CK (n_0_95), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[72][9]  (.Q (\o_values[72] [9] ), .CK (n_0_95), .D (sps__n37));
DFF_X1 \o_values_reg[72][10]  (.Q (\o_values[72] [10] ), .CK (n_0_95), .D (sps__n4));
DFF_X1 \o_values_reg[72][11]  (.Q (\o_values[72] [11] ), .CK (n_0_95), .D (sps__n10));
DFF_X1 \o_values_reg[72][12]  (.Q (\o_values[72] [12] ), .CK (n_0_95), .D (sps__n7));
DFF_X1 \o_values_reg[72][13]  (.Q (\o_values[72] [13] ), .CK (n_0_95), .D (sps__n1));
DFF_X1 \o_values_reg[72][14]  (.Q (\o_values[72] [14] ), .CK (n_0_95), .D (sps__n13));
DFF_X1 \o_values_reg[72][15]  (.Q (\o_values[72] [15] ), .CK (n_0_95), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[72]_reg  (.GCK (n_0_95), .CK (clk), .E (n_0_11), .SE (1'b0 ));
DFF_X1 \o_values_reg[73][0]  (.Q (\o_values[73] [0] ), .CK (n_0_94), .D (sps__n16));
DFF_X1 \o_values_reg[73][1]  (.Q (\o_values[73] [1] ), .CK (n_0_94), .D (sps__n25));
DFF_X1 \o_values_reg[73][2]  (.Q (\o_values[73] [2] ), .CK (n_0_94), .D (sps__n19));
DFF_X1 \o_values_reg[73][3]  (.Q (\o_values[73] [3] ), .CK (n_0_94), .D (sps__n28));
DFF_X1 \o_values_reg[73][4]  (.Q (\o_values[73] [4] ), .CK (n_0_94), .D (sps__n31));
DFF_X1 \o_values_reg[73][5]  (.Q (\o_values[73] [5] ), .CK (n_0_94), .D (sps__n34));
DFF_X1 \o_values_reg[73][6]  (.Q (\o_values[73] [6] ), .CK (n_0_94), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[73][7]  (.Q (\o_values[73] [7] ), .CK (n_0_94), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[73][8]  (.Q (\o_values[73] [8] ), .CK (n_0_94), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[73][9]  (.Q (\o_values[73] [9] ), .CK (n_0_94), .D (sps__n37));
DFF_X1 \o_values_reg[73][10]  (.Q (\o_values[73] [10] ), .CK (n_0_94), .D (sps__n4));
DFF_X1 \o_values_reg[73][11]  (.Q (\o_values[73] [11] ), .CK (n_0_94), .D (sps__n10));
DFF_X1 \o_values_reg[73][12]  (.Q (\o_values[73] [12] ), .CK (n_0_94), .D (sps__n7));
DFF_X1 \o_values_reg[73][13]  (.Q (\o_values[73] [13] ), .CK (n_0_94), .D (sps__n1));
DFF_X1 \o_values_reg[73][14]  (.Q (\o_values[73] [14] ), .CK (n_0_94), .D (sps__n13));
DFF_X1 \o_values_reg[73][15]  (.Q (\o_values[73] [15] ), .CK (n_0_94), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[73]_reg  (.GCK (n_0_94), .CK (clk), .E (n_0_10), .SE (1'b0 ));
DFF_X1 \o_values_reg[74][0]  (.Q (\o_values[74] [0] ), .CK (n_0_93), .D (sps__n16));
DFF_X1 \o_values_reg[74][1]  (.Q (\o_values[74] [1] ), .CK (n_0_93), .D (sps__n25));
DFF_X1 \o_values_reg[74][2]  (.Q (\o_values[74] [2] ), .CK (n_0_93), .D (sps__n19));
DFF_X1 \o_values_reg[74][3]  (.Q (\o_values[74] [3] ), .CK (n_0_93), .D (sps__n28));
DFF_X1 \o_values_reg[74][4]  (.Q (\o_values[74] [4] ), .CK (n_0_93), .D (sps__n31));
DFF_X1 \o_values_reg[74][5]  (.Q (\o_values[74] [5] ), .CK (n_0_93), .D (sps__n34));
DFF_X1 \o_values_reg[74][6]  (.Q (\o_values[74] [6] ), .CK (n_0_93), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[74][7]  (.Q (\o_values[74] [7] ), .CK (n_0_93), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[74][8]  (.Q (\o_values[74] [8] ), .CK (n_0_93), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[74][9]  (.Q (\o_values[74] [9] ), .CK (n_0_93), .D (sps__n37));
DFF_X1 \o_values_reg[74][10]  (.Q (\o_values[74] [10] ), .CK (n_0_93), .D (sps__n4));
DFF_X1 \o_values_reg[74][11]  (.Q (\o_values[74] [11] ), .CK (n_0_93), .D (sps__n10));
DFF_X1 \o_values_reg[74][12]  (.Q (\o_values[74] [12] ), .CK (n_0_93), .D (sps__n7));
DFF_X1 \o_values_reg[74][13]  (.Q (\o_values[74] [13] ), .CK (n_0_93), .D (sps__n1));
DFF_X1 \o_values_reg[74][14]  (.Q (\o_values[74] [14] ), .CK (n_0_93), .D (sps__n13));
DFF_X1 \o_values_reg[74][15]  (.Q (\o_values[74] [15] ), .CK (n_0_93), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[74]_reg  (.GCK (n_0_93), .CK (clk), .E (n_0_9), .SE (1'b0 ));
DFF_X1 \o_values_reg[75][0]  (.Q (\o_values[75] [0] ), .CK (n_0_92), .D (sps__n16));
DFF_X1 \o_values_reg[75][1]  (.Q (\o_values[75] [1] ), .CK (n_0_92), .D (sps__n25));
DFF_X1 \o_values_reg[75][2]  (.Q (\o_values[75] [2] ), .CK (n_0_92), .D (sps__n19));
DFF_X1 \o_values_reg[75][3]  (.Q (\o_values[75] [3] ), .CK (n_0_92), .D (sps__n28));
DFF_X1 \o_values_reg[75][4]  (.Q (\o_values[75] [4] ), .CK (n_0_92), .D (sps__n31));
DFF_X1 \o_values_reg[75][5]  (.Q (\o_values[75] [5] ), .CK (n_0_92), .D (sps__n34));
DFF_X1 \o_values_reg[75][6]  (.Q (\o_values[75] [6] ), .CK (n_0_92), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[75][7]  (.Q (\o_values[75] [7] ), .CK (n_0_92), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[75][8]  (.Q (\o_values[75] [8] ), .CK (n_0_92), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[75][9]  (.Q (\o_values[75] [9] ), .CK (n_0_92), .D (sps__n37));
DFF_X1 \o_values_reg[75][10]  (.Q (\o_values[75] [10] ), .CK (n_0_92), .D (sps__n4));
DFF_X1 \o_values_reg[75][11]  (.Q (\o_values[75] [11] ), .CK (n_0_92), .D (sps__n10));
DFF_X1 \o_values_reg[75][12]  (.Q (\o_values[75] [12] ), .CK (n_0_92), .D (sps__n7));
DFF_X1 \o_values_reg[75][13]  (.Q (\o_values[75] [13] ), .CK (n_0_92), .D (sps__n1));
DFF_X1 \o_values_reg[75][14]  (.Q (\o_values[75] [14] ), .CK (n_0_92), .D (sps__n13));
DFF_X1 \o_values_reg[75][15]  (.Q (\o_values[75] [15] ), .CK (n_0_92), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[75]_reg  (.GCK (n_0_92), .CK (clk), .E (n_0_8), .SE (1'b0 ));
DFF_X1 \o_values_reg[76][0]  (.Q (\o_values[76] [0] ), .CK (n_0_91), .D (sps__n16));
DFF_X1 \o_values_reg[76][1]  (.Q (\o_values[76] [1] ), .CK (n_0_91), .D (sps__n25));
DFF_X1 \o_values_reg[76][2]  (.Q (\o_values[76] [2] ), .CK (n_0_91), .D (sps__n19));
DFF_X1 \o_values_reg[76][3]  (.Q (\o_values[76] [3] ), .CK (n_0_91), .D (sps__n28));
DFF_X1 \o_values_reg[76][4]  (.Q (\o_values[76] [4] ), .CK (n_0_91), .D (sps__n31));
DFF_X1 \o_values_reg[76][5]  (.Q (\o_values[76] [5] ), .CK (n_0_91), .D (sps__n34));
DFF_X1 \o_values_reg[76][6]  (.Q (\o_values[76] [6] ), .CK (n_0_91), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[76][7]  (.Q (\o_values[76] [7] ), .CK (n_0_91), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[76][8]  (.Q (\o_values[76] [8] ), .CK (n_0_91), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[76][9]  (.Q (\o_values[76] [9] ), .CK (n_0_91), .D (sps__n37));
DFF_X1 \o_values_reg[76][10]  (.Q (\o_values[76] [10] ), .CK (n_0_91), .D (sps__n4));
DFF_X1 \o_values_reg[76][11]  (.Q (\o_values[76] [11] ), .CK (n_0_91), .D (sps__n10));
DFF_X1 \o_values_reg[76][12]  (.Q (\o_values[76] [12] ), .CK (n_0_91), .D (sps__n7));
DFF_X1 \o_values_reg[76][13]  (.Q (\o_values[76] [13] ), .CK (n_0_91), .D (sps__n1));
DFF_X1 \o_values_reg[76][14]  (.Q (\o_values[76] [14] ), .CK (n_0_91), .D (sps__n13));
DFF_X1 \o_values_reg[76][15]  (.Q (\o_values[76] [15] ), .CK (n_0_91), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[76]_reg  (.GCK (n_0_91), .CK (clk), .E (n_0_7), .SE (1'b0 ));
DFF_X1 \o_values_reg[77][0]  (.Q (\o_values[77] [0] ), .CK (n_0_90), .D (sps__n16));
DFF_X1 \o_values_reg[77][1]  (.Q (\o_values[77] [1] ), .CK (n_0_90), .D (sps__n25));
DFF_X1 \o_values_reg[77][2]  (.Q (\o_values[77] [2] ), .CK (n_0_90), .D (sps__n19));
DFF_X1 \o_values_reg[77][3]  (.Q (\o_values[77] [3] ), .CK (n_0_90), .D (sps__n28));
DFF_X1 \o_values_reg[77][4]  (.Q (\o_values[77] [4] ), .CK (n_0_90), .D (sps__n31));
DFF_X1 \o_values_reg[77][5]  (.Q (\o_values[77] [5] ), .CK (n_0_90), .D (sps__n34));
DFF_X1 \o_values_reg[77][6]  (.Q (\o_values[77] [6] ), .CK (n_0_90), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[77][7]  (.Q (\o_values[77] [7] ), .CK (n_0_90), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[77][8]  (.Q (\o_values[77] [8] ), .CK (n_0_90), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[77][9]  (.Q (\o_values[77] [9] ), .CK (n_0_90), .D (sps__n37));
DFF_X1 \o_values_reg[77][10]  (.Q (\o_values[77] [10] ), .CK (n_0_90), .D (sps__n4));
DFF_X1 \o_values_reg[77][11]  (.Q (\o_values[77] [11] ), .CK (n_0_90), .D (sps__n10));
DFF_X1 \o_values_reg[77][12]  (.Q (\o_values[77] [12] ), .CK (n_0_90), .D (sps__n7));
DFF_X1 \o_values_reg[77][13]  (.Q (\o_values[77] [13] ), .CK (n_0_90), .D (sps__n1));
DFF_X1 \o_values_reg[77][14]  (.Q (\o_values[77] [14] ), .CK (n_0_90), .D (sps__n13));
DFF_X1 \o_values_reg[77][15]  (.Q (\o_values[77] [15] ), .CK (n_0_90), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[77]_reg  (.GCK (n_0_90), .CK (clk), .E (n_0_6), .SE (1'b0 ));
DFF_X1 \o_values_reg[78][0]  (.Q (\o_values[78] [0] ), .CK (n_0_89), .D (sps__n16));
DFF_X1 \o_values_reg[78][1]  (.Q (\o_values[78] [1] ), .CK (n_0_89), .D (sps__n25));
DFF_X1 \o_values_reg[78][2]  (.Q (\o_values[78] [2] ), .CK (n_0_89), .D (sps__n19));
DFF_X1 \o_values_reg[78][3]  (.Q (\o_values[78] [3] ), .CK (n_0_89), .D (sps__n28));
DFF_X1 \o_values_reg[78][4]  (.Q (\o_values[78] [4] ), .CK (n_0_89), .D (sps__n31));
DFF_X1 \o_values_reg[78][5]  (.Q (\o_values[78] [5] ), .CK (n_0_89), .D (sps__n34));
DFF_X1 \o_values_reg[78][6]  (.Q (\o_values[78] [6] ), .CK (n_0_89), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[78][7]  (.Q (\o_values[78] [7] ), .CK (n_0_89), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[78][8]  (.Q (\o_values[78] [8] ), .CK (n_0_89), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[78][9]  (.Q (\o_values[78] [9] ), .CK (n_0_89), .D (sps__n37));
DFF_X1 \o_values_reg[78][10]  (.Q (\o_values[78] [10] ), .CK (n_0_89), .D (sps__n4));
DFF_X1 \o_values_reg[78][11]  (.Q (\o_values[78] [11] ), .CK (n_0_89), .D (sps__n10));
DFF_X1 \o_values_reg[78][12]  (.Q (\o_values[78] [12] ), .CK (n_0_89), .D (sps__n7));
DFF_X1 \o_values_reg[78][13]  (.Q (\o_values[78] [13] ), .CK (n_0_89), .D (sps__n1));
DFF_X1 \o_values_reg[78][14]  (.Q (\o_values[78] [14] ), .CK (n_0_89), .D (sps__n13));
DFF_X1 \o_values_reg[78][15]  (.Q (\o_values[78] [15] ), .CK (n_0_89), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[78]_reg  (.GCK (n_0_89), .CK (clk), .E (n_0_5), .SE (1'b0 ));
DFF_X1 \o_values_reg[79][0]  (.Q (\o_values[79] [0] ), .CK (n_0_88), .D (sps__n16));
DFF_X1 \o_values_reg[79][1]  (.Q (\o_values[79] [1] ), .CK (n_0_88), .D (sps__n25));
DFF_X1 \o_values_reg[79][2]  (.Q (\o_values[79] [2] ), .CK (n_0_88), .D (sps__n19));
DFF_X1 \o_values_reg[79][3]  (.Q (\o_values[79] [3] ), .CK (n_0_88), .D (sps__n28));
DFF_X1 \o_values_reg[79][4]  (.Q (\o_values[79] [4] ), .CK (n_0_88), .D (sps__n31));
DFF_X1 \o_values_reg[79][5]  (.Q (\o_values[79] [5] ), .CK (n_0_88), .D (sps__n34));
DFF_X1 \o_values_reg[79][6]  (.Q (\o_values[79] [6] ), .CK (n_0_88), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[79][7]  (.Q (\o_values[79] [7] ), .CK (n_0_88), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[79][8]  (.Q (\o_values[79] [8] ), .CK (n_0_88), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[79][9]  (.Q (\o_values[79] [9] ), .CK (n_0_88), .D (sps__n37));
DFF_X1 \o_values_reg[79][10]  (.Q (\o_values[79] [10] ), .CK (n_0_88), .D (sps__n4));
DFF_X1 \o_values_reg[79][11]  (.Q (\o_values[79] [11] ), .CK (n_0_88), .D (sps__n10));
DFF_X1 \o_values_reg[79][12]  (.Q (\o_values[79] [12] ), .CK (n_0_88), .D (sps__n7));
DFF_X1 \o_values_reg[79][13]  (.Q (\o_values[79] [13] ), .CK (n_0_88), .D (sps__n1));
DFF_X1 \o_values_reg[79][14]  (.Q (\o_values[79] [14] ), .CK (n_0_88), .D (sps__n13));
DFF_X1 \o_values_reg[79][15]  (.Q (\o_values[79] [15] ), .CK (n_0_88), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[79]_reg  (.GCK (n_0_88), .CK (clk), .E (n_0_4), .SE (1'b0 ));
DFF_X1 \o_values_reg[80][0]  (.Q (\o_values[80] [0] ), .CK (n_0_87), .D (sps__n16));
DFF_X1 \o_values_reg[80][1]  (.Q (\o_values[80] [1] ), .CK (n_0_87), .D (sps__n25));
DFF_X1 \o_values_reg[80][2]  (.Q (\o_values[80] [2] ), .CK (n_0_87), .D (sps__n19));
DFF_X1 \o_values_reg[80][3]  (.Q (\o_values[80] [3] ), .CK (n_0_87), .D (sps__n28));
DFF_X1 \o_values_reg[80][4]  (.Q (\o_values[80] [4] ), .CK (n_0_87), .D (sps__n31));
DFF_X1 \o_values_reg[80][5]  (.Q (\o_values[80] [5] ), .CK (n_0_87), .D (sps__n34));
DFF_X1 \o_values_reg[80][6]  (.Q (\o_values[80] [6] ), .CK (n_0_87), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[80][7]  (.Q (\o_values[80] [7] ), .CK (n_0_87), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[80][8]  (.Q (\o_values[80] [8] ), .CK (n_0_87), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[80][9]  (.Q (\o_values[80] [9] ), .CK (n_0_87), .D (sps__n37));
DFF_X1 \o_values_reg[80][10]  (.Q (\o_values[80] [10] ), .CK (n_0_87), .D (sps__n4));
DFF_X1 \o_values_reg[80][11]  (.Q (\o_values[80] [11] ), .CK (n_0_87), .D (sps__n10));
DFF_X1 \o_values_reg[80][12]  (.Q (\o_values[80] [12] ), .CK (n_0_87), .D (sps__n7));
DFF_X1 \o_values_reg[80][13]  (.Q (\o_values[80] [13] ), .CK (n_0_87), .D (sps__n1));
DFF_X1 \o_values_reg[80][14]  (.Q (\o_values[80] [14] ), .CK (n_0_87), .D (sps__n13));
DFF_X1 \o_values_reg[80][15]  (.Q (\o_values[80] [15] ), .CK (n_0_87), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[80]_reg  (.GCK (n_0_87), .CK (clk), .E (n_0_3), .SE (1'b0 ));
DFF_X1 \o_values_reg[81][0]  (.Q (\o_values[81] [0] ), .CK (n_0_86), .D (sps__n16));
DFF_X1 \o_values_reg[81][1]  (.Q (\o_values[81] [1] ), .CK (n_0_86), .D (sps__n25));
DFF_X1 \o_values_reg[81][2]  (.Q (\o_values[81] [2] ), .CK (n_0_86), .D (sps__n19));
DFF_X1 \o_values_reg[81][3]  (.Q (\o_values[81] [3] ), .CK (n_0_86), .D (sps__n28));
DFF_X1 \o_values_reg[81][4]  (.Q (\o_values[81] [4] ), .CK (n_0_86), .D (sps__n31));
DFF_X1 \o_values_reg[81][5]  (.Q (\o_values[81] [5] ), .CK (n_0_86), .D (sps__n34));
DFF_X1 \o_values_reg[81][6]  (.Q (\o_values[81] [6] ), .CK (n_0_86), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[81][7]  (.Q (\o_values[81] [7] ), .CK (n_0_86), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[81][8]  (.Q (\o_values[81] [8] ), .CK (n_0_86), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[81][9]  (.Q (\o_values[81] [9] ), .CK (n_0_86), .D (sps__n37));
DFF_X1 \o_values_reg[81][10]  (.Q (\o_values[81] [10] ), .CK (n_0_86), .D (sps__n4));
DFF_X1 \o_values_reg[81][11]  (.Q (\o_values[81] [11] ), .CK (n_0_86), .D (sps__n10));
DFF_X1 \o_values_reg[81][12]  (.Q (\o_values[81] [12] ), .CK (n_0_86), .D (sps__n7));
DFF_X1 \o_values_reg[81][13]  (.Q (\o_values[81] [13] ), .CK (n_0_86), .D (sps__n1));
DFF_X1 \o_values_reg[81][14]  (.Q (\o_values[81] [14] ), .CK (n_0_86), .D (sps__n13));
DFF_X1 \o_values_reg[81][15]  (.Q (\o_values[81] [15] ), .CK (n_0_86), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[81]_reg  (.GCK (n_0_86), .CK (clk), .E (n_0_2), .SE (1'b0 ));
DFF_X1 \o_values_reg[82][0]  (.Q (\o_values[82] [0] ), .CK (n_0_85), .D (sps__n16));
DFF_X1 \o_values_reg[82][1]  (.Q (\o_values[82] [1] ), .CK (n_0_85), .D (sps__n25));
DFF_X1 \o_values_reg[82][2]  (.Q (\o_values[82] [2] ), .CK (n_0_85), .D (sps__n19));
DFF_X1 \o_values_reg[82][3]  (.Q (\o_values[82] [3] ), .CK (n_0_85), .D (sps__n28));
DFF_X1 \o_values_reg[82][4]  (.Q (\o_values[82] [4] ), .CK (n_0_85), .D (sps__n31));
DFF_X1 \o_values_reg[82][5]  (.Q (\o_values[82] [5] ), .CK (n_0_85), .D (sps__n34));
DFF_X1 \o_values_reg[82][6]  (.Q (\o_values[82] [6] ), .CK (n_0_85), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[82][7]  (.Q (\o_values[82] [7] ), .CK (n_0_85), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[82][8]  (.Q (\o_values[82] [8] ), .CK (n_0_85), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[82][9]  (.Q (\o_values[82] [9] ), .CK (n_0_85), .D (sps__n37));
DFF_X1 \o_values_reg[82][10]  (.Q (\o_values[82] [10] ), .CK (n_0_85), .D (sps__n4));
DFF_X1 \o_values_reg[82][11]  (.Q (\o_values[82] [11] ), .CK (n_0_85), .D (sps__n10));
DFF_X1 \o_values_reg[82][12]  (.Q (\o_values[82] [12] ), .CK (n_0_85), .D (sps__n7));
DFF_X1 \o_values_reg[82][13]  (.Q (\o_values[82] [13] ), .CK (n_0_85), .D (sps__n1));
DFF_X1 \o_values_reg[82][14]  (.Q (\o_values[82] [14] ), .CK (n_0_85), .D (sps__n13));
DFF_X1 \o_values_reg[82][15]  (.Q (\o_values[82] [15] ), .CK (n_0_85), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[82]_reg  (.GCK (n_0_85), .CK (clk), .E (n_0_1), .SE (1'b0 ));
DFF_X1 \o_values_reg[83][0]  (.Q (\o_values[83] [0] ), .CK (n_0_84), .D (sps__n16));
DFF_X1 \o_values_reg[83][1]  (.Q (\o_values[83] [1] ), .CK (n_0_84), .D (sps__n25));
DFF_X1 \o_values_reg[83][2]  (.Q (\o_values[83] [2] ), .CK (n_0_84), .D (sps__n19));
DFF_X1 \o_values_reg[83][3]  (.Q (\o_values[83] [3] ), .CK (n_0_84), .D (sps__n28));
DFF_X1 \o_values_reg[83][4]  (.Q (\o_values[83] [4] ), .CK (n_0_84), .D (sps__n31));
DFF_X1 \o_values_reg[83][5]  (.Q (\o_values[83] [5] ), .CK (n_0_84), .D (sps__n34));
DFF_X1 \o_values_reg[83][6]  (.Q (\o_values[83] [6] ), .CK (n_0_84), .D (\t_o_values[6] ));
DFF_X1 \o_values_reg[83][7]  (.Q (\o_values[83] [7] ), .CK (n_0_84), .D (\t_o_values[7] ));
DFF_X1 \o_values_reg[83][8]  (.Q (\o_values[83] [8] ), .CK (n_0_84), .D (\t_o_values[8] ));
DFF_X1 \o_values_reg[83][9]  (.Q (\o_values[83] [9] ), .CK (n_0_84), .D (sps__n37));
DFF_X1 \o_values_reg[83][10]  (.Q (\o_values[83] [10] ), .CK (n_0_84), .D (sps__n4));
DFF_X1 \o_values_reg[83][11]  (.Q (\o_values[83] [11] ), .CK (n_0_84), .D (sps__n10));
DFF_X1 \o_values_reg[83][12]  (.Q (\o_values[83] [12] ), .CK (n_0_84), .D (sps__n7));
DFF_X1 \o_values_reg[83][13]  (.Q (\o_values[83] [13] ), .CK (n_0_84), .D (sps__n1));
DFF_X1 \o_values_reg[83][14]  (.Q (\o_values[83] [14] ), .CK (n_0_84), .D (sps__n13));
DFF_X1 \o_values_reg[83][15]  (.Q (\o_values[83] [15] ), .CK (n_0_84), .D (sps__n22));
CLKGATETST_X1 \clk_gate_o_values_reg[83]_reg  (.GCK (n_0_84), .CK (clk), .E (n_0_0), .SE (1'b0 ));
BUF_X8 sps__L1_c1 (.Z (sps__n1), .A (\t_o_values[13] ));
BUF_X8 sps__L1_c4 (.Z (sps__n4), .A (\t_o_values[10] ));
BUF_X8 sps__L1_c7 (.Z (sps__n7), .A (\t_o_values[12] ));
BUF_X8 sps__L1_c10 (.Z (sps__n10), .A (\t_o_values[11] ));
BUF_X8 sps__L1_c13 (.Z (sps__n13), .A (\t_o_values[14] ));
BUF_X8 sps__L1_c16 (.Z (sps__n16), .A (\t_o_values[0] ));
BUF_X8 sps__L1_c19 (.Z (sps__n19), .A (\t_o_values[2] ));
BUF_X8 sps__L1_c22 (.Z (sps__n22), .A (\t_o_values[15] ));
BUF_X8 sps__L1_c25 (.Z (sps__n25), .A (\t_o_values[1] ));
BUF_X8 sps__L1_c28 (.Z (sps__n28), .A (\t_o_values[3] ));
BUF_X8 sps__L1_c31 (.Z (sps__n31), .A (\t_o_values[4] ));
BUF_X8 sps__L1_c34 (.Z (sps__n34), .A (\t_o_values[5] ));
BUF_X8 sps__L1_c37 (.Z (sps__n37), .A (\t_o_values[9] ));

endmodule //Neuron_Layer


