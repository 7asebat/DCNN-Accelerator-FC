/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 23:27:34 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3521584009 */

module Neuron_Layer(clk, load_en, load_value, load_address, reset, \o_values[0] , 
      \o_values[1] , \o_values[2] , \o_values[3] , \o_values[4] , \o_values[5] , 
      \o_values[6] , \o_values[7] , \o_values[8] , \o_values[9] , \o_values[10] , 
      \o_values[11] , \o_values[12] , \o_values[13] , \o_values[14] , 
      \o_values[15] , \o_values[16] , \o_values[17] , \o_values[18] , 
      \o_values[19] , \o_values[20] , \o_values[21] , \o_values[22] , 
      \o_values[23] , \o_values[24] , \o_values[25] , \o_values[26] , 
      \o_values[27] , \o_values[28] , \o_values[29] , \o_values[30] , 
      \o_values[31] , \o_values[32] , \o_values[33] , \o_values[34] , 
      \o_values[35] , \o_values[36] , \o_values[37] , \o_values[38] , 
      \o_values[39] , \o_values[40] , \o_values[41] , \o_values[42] , 
      \o_values[43] , \o_values[44] , \o_values[45] , \o_values[46] , 
      \o_values[47] , \o_values[48] , \o_values[49] , \o_values[50] , 
      \o_values[51] , \o_values[52] , \o_values[53] , \o_values[54] , 
      \o_values[55] , \o_values[56] , \o_values[57] , \o_values[58] , 
      \o_values[59] , \o_values[60] , \o_values[61] , \o_values[62] , 
      \o_values[63] , \o_values[64] , \o_values[65] , \o_values[66] , 
      \o_values[67] , \o_values[68] , \o_values[69] , \o_values[70] , 
      \o_values[71] , \o_values[72] , \o_values[73] , \o_values[74] , 
      \o_values[75] , \o_values[76] , \o_values[77] , \o_values[78] , 
      \o_values[79] , \o_values[80] , \o_values[81] , \o_values[82] , 
      \o_values[83] );
   input clk;
   input load_en;
   input [15:0]load_value;
   input [15:0]load_address;
   input reset;
   output [15:0]\o_values[0] ;
   output [15:0]\o_values[1] ;
   output [15:0]\o_values[2] ;
   output [15:0]\o_values[3] ;
   output [15:0]\o_values[4] ;
   output [15:0]\o_values[5] ;
   output [15:0]\o_values[6] ;
   output [15:0]\o_values[7] ;
   output [15:0]\o_values[8] ;
   output [15:0]\o_values[9] ;
   output [15:0]\o_values[10] ;
   output [15:0]\o_values[11] ;
   output [15:0]\o_values[12] ;
   output [15:0]\o_values[13] ;
   output [15:0]\o_values[14] ;
   output [15:0]\o_values[15] ;
   output [15:0]\o_values[16] ;
   output [15:0]\o_values[17] ;
   output [15:0]\o_values[18] ;
   output [15:0]\o_values[19] ;
   output [15:0]\o_values[20] ;
   output [15:0]\o_values[21] ;
   output [15:0]\o_values[22] ;
   output [15:0]\o_values[23] ;
   output [15:0]\o_values[24] ;
   output [15:0]\o_values[25] ;
   output [15:0]\o_values[26] ;
   output [15:0]\o_values[27] ;
   output [15:0]\o_values[28] ;
   output [15:0]\o_values[29] ;
   output [15:0]\o_values[30] ;
   output [15:0]\o_values[31] ;
   output [15:0]\o_values[32] ;
   output [15:0]\o_values[33] ;
   output [15:0]\o_values[34] ;
   output [15:0]\o_values[35] ;
   output [15:0]\o_values[36] ;
   output [15:0]\o_values[37] ;
   output [15:0]\o_values[38] ;
   output [15:0]\o_values[39] ;
   output [15:0]\o_values[40] ;
   output [15:0]\o_values[41] ;
   output [15:0]\o_values[42] ;
   output [15:0]\o_values[43] ;
   output [15:0]\o_values[44] ;
   output [15:0]\o_values[45] ;
   output [15:0]\o_values[46] ;
   output [15:0]\o_values[47] ;
   output [15:0]\o_values[48] ;
   output [15:0]\o_values[49] ;
   output [15:0]\o_values[50] ;
   output [15:0]\o_values[51] ;
   output [15:0]\o_values[52] ;
   output [15:0]\o_values[53] ;
   output [15:0]\o_values[54] ;
   output [15:0]\o_values[55] ;
   output [15:0]\o_values[56] ;
   output [15:0]\o_values[57] ;
   output [15:0]\o_values[58] ;
   output [15:0]\o_values[59] ;
   output [15:0]\o_values[60] ;
   output [15:0]\o_values[61] ;
   output [15:0]\o_values[62] ;
   output [15:0]\o_values[63] ;
   output [15:0]\o_values[64] ;
   output [15:0]\o_values[65] ;
   output [15:0]\o_values[66] ;
   output [15:0]\o_values[67] ;
   output [15:0]\o_values[68] ;
   output [15:0]\o_values[69] ;
   output [15:0]\o_values[70] ;
   output [15:0]\o_values[71] ;
   output [15:0]\o_values[72] ;
   output [15:0]\o_values[73] ;
   output [15:0]\o_values[74] ;
   output [15:0]\o_values[75] ;
   output [15:0]\o_values[76] ;
   output [15:0]\o_values[77] ;
   output [15:0]\o_values[78] ;
   output [15:0]\o_values[79] ;
   output [15:0]\o_values[80] ;
   output [15:0]\o_values[81] ;
   output [15:0]\o_values[82] ;
   output [15:0]\o_values[83] ;

   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire [15:0]o_values;
   wire n_0_83;
   wire n_0_82;
   wire n_0_81;
   wire n_0_80;
   wire n_0_0_0;
   wire n_0_79;
   wire n_0_78;
   wire n_0_77;
   wire n_0_76;
   wire n_0_0_1;
   wire n_0_75;
   wire n_0_74;
   wire n_0_73;
   wire n_0_72;
   wire n_0_0_2;
   wire n_0_71;
   wire n_0_70;
   wire n_0_69;
   wire n_0_68;
   wire n_0_0_3;
   wire n_0_67;
   wire n_0_66;
   wire n_0_65;
   wire n_0_64;
   wire n_0_63;
   wire n_0_62;
   wire n_0_61;
   wire n_0_60;
   wire n_0_0_4;
   wire n_0_59;
   wire n_0_58;
   wire n_0_57;
   wire n_0_56;
   wire n_0_0_5;
   wire n_0_55;
   wire n_0_54;
   wire n_0_53;
   wire n_0_52;
   wire n_0_0_6;
   wire n_0_51;
   wire n_0_50;
   wire n_0_49;
   wire n_0_48;
   wire n_0_0_7;
   wire n_0_47;
   wire n_0_46;
   wire n_0_45;
   wire n_0_44;
   wire n_0_0_8;
   wire n_0_43;
   wire n_0_42;
   wire n_0_41;
   wire n_0_40;
   wire n_0_0_9;
   wire n_0_39;
   wire n_0_38;
   wire n_0_37;
   wire n_0_36;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_35;
   wire n_0_34;
   wire n_0_33;
   wire n_0_32;
   wire n_0_0_12;
   wire n_0_31;
   wire n_0_30;
   wire n_0_29;
   wire n_0_28;
   wire n_0_0_13;
   wire n_0_27;
   wire n_0_26;
   wire n_0_25;
   wire n_0_24;
   wire n_0_0_14;
   wire n_0_23;
   wire n_0_0_15;
   wire n_0_22;
   wire n_0_0_16;
   wire n_0_21;
   wire n_0_0_17;
   wire n_0_20;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_19;
   wire n_0_18;
   wire n_0_17;
   wire n_0_16;
   wire n_0_15;
   wire n_0_14;
   wire n_0_13;
   wire n_0_12;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_11;
   wire n_0_10;
   wire n_0_9;
   wire n_0_8;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_7;
   wire n_0_0_25;
   wire n_0_6;
   wire n_0_0_26;
   wire n_0_5;
   wire n_0_0_27;
   wire n_0_4;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_3;
   wire n_0_0_33;
   wire n_0_2;
   wire n_0_0_34;
   wire n_0_1;
   wire n_0_0_35;
   wire n_0_0;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;

   CLKGATETST_X1 \clk_gate_o_values_reg[83]_reg  (.CK(clk), .E(n_0_0), .SE(1'b0), 
      .GCK(n_0_84));
   DFF_X1 \o_values_reg[83][15]  (.D(o_values[15]), .CK(n_0_84), .Q(
      \o_values[83] [15]), .QN());
   DFF_X1 \o_values_reg[83][14]  (.D(o_values[14]), .CK(n_0_84), .Q(
      \o_values[83] [14]), .QN());
   DFF_X1 \o_values_reg[83][13]  (.D(o_values[13]), .CK(n_0_84), .Q(
      \o_values[83] [13]), .QN());
   DFF_X1 \o_values_reg[83][12]  (.D(o_values[12]), .CK(n_0_84), .Q(
      \o_values[83] [12]), .QN());
   DFF_X1 \o_values_reg[83][11]  (.D(o_values[11]), .CK(n_0_84), .Q(
      \o_values[83] [11]), .QN());
   DFF_X1 \o_values_reg[83][10]  (.D(o_values[10]), .CK(n_0_84), .Q(
      \o_values[83] [10]), .QN());
   DFF_X1 \o_values_reg[83][9]  (.D(o_values[9]), .CK(n_0_84), .Q(
      \o_values[83] [9]), .QN());
   DFF_X1 \o_values_reg[83][8]  (.D(o_values[8]), .CK(n_0_84), .Q(
      \o_values[83] [8]), .QN());
   DFF_X1 \o_values_reg[83][7]  (.D(o_values[7]), .CK(n_0_84), .Q(
      \o_values[83] [7]), .QN());
   DFF_X1 \o_values_reg[83][6]  (.D(o_values[6]), .CK(n_0_84), .Q(
      \o_values[83] [6]), .QN());
   DFF_X1 \o_values_reg[83][5]  (.D(o_values[5]), .CK(n_0_84), .Q(
      \o_values[83] [5]), .QN());
   DFF_X1 \o_values_reg[83][4]  (.D(o_values[4]), .CK(n_0_84), .Q(
      \o_values[83] [4]), .QN());
   DFF_X1 \o_values_reg[83][3]  (.D(o_values[3]), .CK(n_0_84), .Q(
      \o_values[83] [3]), .QN());
   DFF_X1 \o_values_reg[83][2]  (.D(o_values[2]), .CK(n_0_84), .Q(
      \o_values[83] [2]), .QN());
   DFF_X1 \o_values_reg[83][1]  (.D(o_values[1]), .CK(n_0_84), .Q(
      \o_values[83] [1]), .QN());
   DFF_X1 \o_values_reg[83][0]  (.D(o_values[0]), .CK(n_0_84), .Q(
      \o_values[83] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[82]_reg  (.CK(clk), .E(n_0_1), .SE(1'b0), 
      .GCK(n_0_85));
   DFF_X1 \o_values_reg[82][15]  (.D(o_values[15]), .CK(n_0_85), .Q(
      \o_values[82] [15]), .QN());
   DFF_X1 \o_values_reg[82][14]  (.D(o_values[14]), .CK(n_0_85), .Q(
      \o_values[82] [14]), .QN());
   DFF_X1 \o_values_reg[82][13]  (.D(o_values[13]), .CK(n_0_85), .Q(
      \o_values[82] [13]), .QN());
   DFF_X1 \o_values_reg[82][12]  (.D(o_values[12]), .CK(n_0_85), .Q(
      \o_values[82] [12]), .QN());
   DFF_X1 \o_values_reg[82][11]  (.D(o_values[11]), .CK(n_0_85), .Q(
      \o_values[82] [11]), .QN());
   DFF_X1 \o_values_reg[82][10]  (.D(o_values[10]), .CK(n_0_85), .Q(
      \o_values[82] [10]), .QN());
   DFF_X1 \o_values_reg[82][9]  (.D(o_values[9]), .CK(n_0_85), .Q(
      \o_values[82] [9]), .QN());
   DFF_X1 \o_values_reg[82][8]  (.D(o_values[8]), .CK(n_0_85), .Q(
      \o_values[82] [8]), .QN());
   DFF_X1 \o_values_reg[82][7]  (.D(o_values[7]), .CK(n_0_85), .Q(
      \o_values[82] [7]), .QN());
   DFF_X1 \o_values_reg[82][6]  (.D(o_values[6]), .CK(n_0_85), .Q(
      \o_values[82] [6]), .QN());
   DFF_X1 \o_values_reg[82][5]  (.D(o_values[5]), .CK(n_0_85), .Q(
      \o_values[82] [5]), .QN());
   DFF_X1 \o_values_reg[82][4]  (.D(o_values[4]), .CK(n_0_85), .Q(
      \o_values[82] [4]), .QN());
   DFF_X1 \o_values_reg[82][3]  (.D(o_values[3]), .CK(n_0_85), .Q(
      \o_values[82] [3]), .QN());
   DFF_X1 \o_values_reg[82][2]  (.D(o_values[2]), .CK(n_0_85), .Q(
      \o_values[82] [2]), .QN());
   DFF_X1 \o_values_reg[82][1]  (.D(o_values[1]), .CK(n_0_85), .Q(
      \o_values[82] [1]), .QN());
   DFF_X1 \o_values_reg[82][0]  (.D(o_values[0]), .CK(n_0_85), .Q(
      \o_values[82] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[81]_reg  (.CK(clk), .E(n_0_2), .SE(1'b0), 
      .GCK(n_0_86));
   DFF_X1 \o_values_reg[81][15]  (.D(o_values[15]), .CK(n_0_86), .Q(
      \o_values[81] [15]), .QN());
   DFF_X1 \o_values_reg[81][14]  (.D(o_values[14]), .CK(n_0_86), .Q(
      \o_values[81] [14]), .QN());
   DFF_X1 \o_values_reg[81][13]  (.D(o_values[13]), .CK(n_0_86), .Q(
      \o_values[81] [13]), .QN());
   DFF_X1 \o_values_reg[81][12]  (.D(o_values[12]), .CK(n_0_86), .Q(
      \o_values[81] [12]), .QN());
   DFF_X1 \o_values_reg[81][11]  (.D(o_values[11]), .CK(n_0_86), .Q(
      \o_values[81] [11]), .QN());
   DFF_X1 \o_values_reg[81][10]  (.D(o_values[10]), .CK(n_0_86), .Q(
      \o_values[81] [10]), .QN());
   DFF_X1 \o_values_reg[81][9]  (.D(o_values[9]), .CK(n_0_86), .Q(
      \o_values[81] [9]), .QN());
   DFF_X1 \o_values_reg[81][8]  (.D(o_values[8]), .CK(n_0_86), .Q(
      \o_values[81] [8]), .QN());
   DFF_X1 \o_values_reg[81][7]  (.D(o_values[7]), .CK(n_0_86), .Q(
      \o_values[81] [7]), .QN());
   DFF_X1 \o_values_reg[81][6]  (.D(o_values[6]), .CK(n_0_86), .Q(
      \o_values[81] [6]), .QN());
   DFF_X1 \o_values_reg[81][5]  (.D(o_values[5]), .CK(n_0_86), .Q(
      \o_values[81] [5]), .QN());
   DFF_X1 \o_values_reg[81][4]  (.D(o_values[4]), .CK(n_0_86), .Q(
      \o_values[81] [4]), .QN());
   DFF_X1 \o_values_reg[81][3]  (.D(o_values[3]), .CK(n_0_86), .Q(
      \o_values[81] [3]), .QN());
   DFF_X1 \o_values_reg[81][2]  (.D(o_values[2]), .CK(n_0_86), .Q(
      \o_values[81] [2]), .QN());
   DFF_X1 \o_values_reg[81][1]  (.D(o_values[1]), .CK(n_0_86), .Q(
      \o_values[81] [1]), .QN());
   DFF_X1 \o_values_reg[81][0]  (.D(o_values[0]), .CK(n_0_86), .Q(
      \o_values[81] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[80]_reg  (.CK(clk), .E(n_0_3), .SE(1'b0), 
      .GCK(n_0_87));
   DFF_X1 \o_values_reg[80][15]  (.D(o_values[15]), .CK(n_0_87), .Q(
      \o_values[80] [15]), .QN());
   DFF_X1 \o_values_reg[80][14]  (.D(o_values[14]), .CK(n_0_87), .Q(
      \o_values[80] [14]), .QN());
   DFF_X1 \o_values_reg[80][13]  (.D(o_values[13]), .CK(n_0_87), .Q(
      \o_values[80] [13]), .QN());
   DFF_X1 \o_values_reg[80][12]  (.D(o_values[12]), .CK(n_0_87), .Q(
      \o_values[80] [12]), .QN());
   DFF_X1 \o_values_reg[80][11]  (.D(o_values[11]), .CK(n_0_87), .Q(
      \o_values[80] [11]), .QN());
   DFF_X1 \o_values_reg[80][10]  (.D(o_values[10]), .CK(n_0_87), .Q(
      \o_values[80] [10]), .QN());
   DFF_X1 \o_values_reg[80][9]  (.D(o_values[9]), .CK(n_0_87), .Q(
      \o_values[80] [9]), .QN());
   DFF_X1 \o_values_reg[80][8]  (.D(o_values[8]), .CK(n_0_87), .Q(
      \o_values[80] [8]), .QN());
   DFF_X1 \o_values_reg[80][7]  (.D(o_values[7]), .CK(n_0_87), .Q(
      \o_values[80] [7]), .QN());
   DFF_X1 \o_values_reg[80][6]  (.D(o_values[6]), .CK(n_0_87), .Q(
      \o_values[80] [6]), .QN());
   DFF_X1 \o_values_reg[80][5]  (.D(o_values[5]), .CK(n_0_87), .Q(
      \o_values[80] [5]), .QN());
   DFF_X1 \o_values_reg[80][4]  (.D(o_values[4]), .CK(n_0_87), .Q(
      \o_values[80] [4]), .QN());
   DFF_X1 \o_values_reg[80][3]  (.D(o_values[3]), .CK(n_0_87), .Q(
      \o_values[80] [3]), .QN());
   DFF_X1 \o_values_reg[80][2]  (.D(o_values[2]), .CK(n_0_87), .Q(
      \o_values[80] [2]), .QN());
   DFF_X1 \o_values_reg[80][1]  (.D(o_values[1]), .CK(n_0_87), .Q(
      \o_values[80] [1]), .QN());
   DFF_X1 \o_values_reg[80][0]  (.D(o_values[0]), .CK(n_0_87), .Q(
      \o_values[80] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[79]_reg  (.CK(clk), .E(n_0_4), .SE(1'b0), 
      .GCK(n_0_88));
   DFF_X1 \o_values_reg[79][15]  (.D(o_values[15]), .CK(n_0_88), .Q(
      \o_values[79] [15]), .QN());
   DFF_X1 \o_values_reg[79][14]  (.D(o_values[14]), .CK(n_0_88), .Q(
      \o_values[79] [14]), .QN());
   DFF_X1 \o_values_reg[79][13]  (.D(o_values[13]), .CK(n_0_88), .Q(
      \o_values[79] [13]), .QN());
   DFF_X1 \o_values_reg[79][12]  (.D(o_values[12]), .CK(n_0_88), .Q(
      \o_values[79] [12]), .QN());
   DFF_X1 \o_values_reg[79][11]  (.D(o_values[11]), .CK(n_0_88), .Q(
      \o_values[79] [11]), .QN());
   DFF_X1 \o_values_reg[79][10]  (.D(o_values[10]), .CK(n_0_88), .Q(
      \o_values[79] [10]), .QN());
   DFF_X1 \o_values_reg[79][9]  (.D(o_values[9]), .CK(n_0_88), .Q(
      \o_values[79] [9]), .QN());
   DFF_X1 \o_values_reg[79][8]  (.D(o_values[8]), .CK(n_0_88), .Q(
      \o_values[79] [8]), .QN());
   DFF_X1 \o_values_reg[79][7]  (.D(o_values[7]), .CK(n_0_88), .Q(
      \o_values[79] [7]), .QN());
   DFF_X1 \o_values_reg[79][6]  (.D(o_values[6]), .CK(n_0_88), .Q(
      \o_values[79] [6]), .QN());
   DFF_X1 \o_values_reg[79][5]  (.D(o_values[5]), .CK(n_0_88), .Q(
      \o_values[79] [5]), .QN());
   DFF_X1 \o_values_reg[79][4]  (.D(o_values[4]), .CK(n_0_88), .Q(
      \o_values[79] [4]), .QN());
   DFF_X1 \o_values_reg[79][3]  (.D(o_values[3]), .CK(n_0_88), .Q(
      \o_values[79] [3]), .QN());
   DFF_X1 \o_values_reg[79][2]  (.D(o_values[2]), .CK(n_0_88), .Q(
      \o_values[79] [2]), .QN());
   DFF_X1 \o_values_reg[79][1]  (.D(o_values[1]), .CK(n_0_88), .Q(
      \o_values[79] [1]), .QN());
   DFF_X1 \o_values_reg[79][0]  (.D(o_values[0]), .CK(n_0_88), .Q(
      \o_values[79] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[78]_reg  (.CK(clk), .E(n_0_5), .SE(1'b0), 
      .GCK(n_0_89));
   DFF_X1 \o_values_reg[78][15]  (.D(o_values[15]), .CK(n_0_89), .Q(
      \o_values[78] [15]), .QN());
   DFF_X1 \o_values_reg[78][14]  (.D(o_values[14]), .CK(n_0_89), .Q(
      \o_values[78] [14]), .QN());
   DFF_X1 \o_values_reg[78][13]  (.D(o_values[13]), .CK(n_0_89), .Q(
      \o_values[78] [13]), .QN());
   DFF_X1 \o_values_reg[78][12]  (.D(o_values[12]), .CK(n_0_89), .Q(
      \o_values[78] [12]), .QN());
   DFF_X1 \o_values_reg[78][11]  (.D(o_values[11]), .CK(n_0_89), .Q(
      \o_values[78] [11]), .QN());
   DFF_X1 \o_values_reg[78][10]  (.D(o_values[10]), .CK(n_0_89), .Q(
      \o_values[78] [10]), .QN());
   DFF_X1 \o_values_reg[78][9]  (.D(o_values[9]), .CK(n_0_89), .Q(
      \o_values[78] [9]), .QN());
   DFF_X1 \o_values_reg[78][8]  (.D(o_values[8]), .CK(n_0_89), .Q(
      \o_values[78] [8]), .QN());
   DFF_X1 \o_values_reg[78][7]  (.D(o_values[7]), .CK(n_0_89), .Q(
      \o_values[78] [7]), .QN());
   DFF_X1 \o_values_reg[78][6]  (.D(o_values[6]), .CK(n_0_89), .Q(
      \o_values[78] [6]), .QN());
   DFF_X1 \o_values_reg[78][5]  (.D(o_values[5]), .CK(n_0_89), .Q(
      \o_values[78] [5]), .QN());
   DFF_X1 \o_values_reg[78][4]  (.D(o_values[4]), .CK(n_0_89), .Q(
      \o_values[78] [4]), .QN());
   DFF_X1 \o_values_reg[78][3]  (.D(o_values[3]), .CK(n_0_89), .Q(
      \o_values[78] [3]), .QN());
   DFF_X1 \o_values_reg[78][2]  (.D(o_values[2]), .CK(n_0_89), .Q(
      \o_values[78] [2]), .QN());
   DFF_X1 \o_values_reg[78][1]  (.D(o_values[1]), .CK(n_0_89), .Q(
      \o_values[78] [1]), .QN());
   DFF_X1 \o_values_reg[78][0]  (.D(o_values[0]), .CK(n_0_89), .Q(
      \o_values[78] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[77]_reg  (.CK(clk), .E(n_0_6), .SE(1'b0), 
      .GCK(n_0_90));
   DFF_X1 \o_values_reg[77][15]  (.D(o_values[15]), .CK(n_0_90), .Q(
      \o_values[77] [15]), .QN());
   DFF_X1 \o_values_reg[77][14]  (.D(o_values[14]), .CK(n_0_90), .Q(
      \o_values[77] [14]), .QN());
   DFF_X1 \o_values_reg[77][13]  (.D(o_values[13]), .CK(n_0_90), .Q(
      \o_values[77] [13]), .QN());
   DFF_X1 \o_values_reg[77][12]  (.D(o_values[12]), .CK(n_0_90), .Q(
      \o_values[77] [12]), .QN());
   DFF_X1 \o_values_reg[77][11]  (.D(o_values[11]), .CK(n_0_90), .Q(
      \o_values[77] [11]), .QN());
   DFF_X1 \o_values_reg[77][10]  (.D(o_values[10]), .CK(n_0_90), .Q(
      \o_values[77] [10]), .QN());
   DFF_X1 \o_values_reg[77][9]  (.D(o_values[9]), .CK(n_0_90), .Q(
      \o_values[77] [9]), .QN());
   DFF_X1 \o_values_reg[77][8]  (.D(o_values[8]), .CK(n_0_90), .Q(
      \o_values[77] [8]), .QN());
   DFF_X1 \o_values_reg[77][7]  (.D(o_values[7]), .CK(n_0_90), .Q(
      \o_values[77] [7]), .QN());
   DFF_X1 \o_values_reg[77][6]  (.D(o_values[6]), .CK(n_0_90), .Q(
      \o_values[77] [6]), .QN());
   DFF_X1 \o_values_reg[77][5]  (.D(o_values[5]), .CK(n_0_90), .Q(
      \o_values[77] [5]), .QN());
   DFF_X1 \o_values_reg[77][4]  (.D(o_values[4]), .CK(n_0_90), .Q(
      \o_values[77] [4]), .QN());
   DFF_X1 \o_values_reg[77][3]  (.D(o_values[3]), .CK(n_0_90), .Q(
      \o_values[77] [3]), .QN());
   DFF_X1 \o_values_reg[77][2]  (.D(o_values[2]), .CK(n_0_90), .Q(
      \o_values[77] [2]), .QN());
   DFF_X1 \o_values_reg[77][1]  (.D(o_values[1]), .CK(n_0_90), .Q(
      \o_values[77] [1]), .QN());
   DFF_X1 \o_values_reg[77][0]  (.D(o_values[0]), .CK(n_0_90), .Q(
      \o_values[77] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[76]_reg  (.CK(clk), .E(n_0_7), .SE(1'b0), 
      .GCK(n_0_91));
   DFF_X1 \o_values_reg[76][15]  (.D(o_values[15]), .CK(n_0_91), .Q(
      \o_values[76] [15]), .QN());
   DFF_X1 \o_values_reg[76][14]  (.D(o_values[14]), .CK(n_0_91), .Q(
      \o_values[76] [14]), .QN());
   DFF_X1 \o_values_reg[76][13]  (.D(o_values[13]), .CK(n_0_91), .Q(
      \o_values[76] [13]), .QN());
   DFF_X1 \o_values_reg[76][12]  (.D(o_values[12]), .CK(n_0_91), .Q(
      \o_values[76] [12]), .QN());
   DFF_X1 \o_values_reg[76][11]  (.D(o_values[11]), .CK(n_0_91), .Q(
      \o_values[76] [11]), .QN());
   DFF_X1 \o_values_reg[76][10]  (.D(o_values[10]), .CK(n_0_91), .Q(
      \o_values[76] [10]), .QN());
   DFF_X1 \o_values_reg[76][9]  (.D(o_values[9]), .CK(n_0_91), .Q(
      \o_values[76] [9]), .QN());
   DFF_X1 \o_values_reg[76][8]  (.D(o_values[8]), .CK(n_0_91), .Q(
      \o_values[76] [8]), .QN());
   DFF_X1 \o_values_reg[76][7]  (.D(o_values[7]), .CK(n_0_91), .Q(
      \o_values[76] [7]), .QN());
   DFF_X1 \o_values_reg[76][6]  (.D(o_values[6]), .CK(n_0_91), .Q(
      \o_values[76] [6]), .QN());
   DFF_X1 \o_values_reg[76][5]  (.D(o_values[5]), .CK(n_0_91), .Q(
      \o_values[76] [5]), .QN());
   DFF_X1 \o_values_reg[76][4]  (.D(o_values[4]), .CK(n_0_91), .Q(
      \o_values[76] [4]), .QN());
   DFF_X1 \o_values_reg[76][3]  (.D(o_values[3]), .CK(n_0_91), .Q(
      \o_values[76] [3]), .QN());
   DFF_X1 \o_values_reg[76][2]  (.D(o_values[2]), .CK(n_0_91), .Q(
      \o_values[76] [2]), .QN());
   DFF_X1 \o_values_reg[76][1]  (.D(o_values[1]), .CK(n_0_91), .Q(
      \o_values[76] [1]), .QN());
   DFF_X1 \o_values_reg[76][0]  (.D(o_values[0]), .CK(n_0_91), .Q(
      \o_values[76] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[75]_reg  (.CK(clk), .E(n_0_8), .SE(1'b0), 
      .GCK(n_0_92));
   DFF_X1 \o_values_reg[75][15]  (.D(o_values[15]), .CK(n_0_92), .Q(
      \o_values[75] [15]), .QN());
   DFF_X1 \o_values_reg[75][14]  (.D(o_values[14]), .CK(n_0_92), .Q(
      \o_values[75] [14]), .QN());
   DFF_X1 \o_values_reg[75][13]  (.D(o_values[13]), .CK(n_0_92), .Q(
      \o_values[75] [13]), .QN());
   DFF_X1 \o_values_reg[75][12]  (.D(o_values[12]), .CK(n_0_92), .Q(
      \o_values[75] [12]), .QN());
   DFF_X1 \o_values_reg[75][11]  (.D(o_values[11]), .CK(n_0_92), .Q(
      \o_values[75] [11]), .QN());
   DFF_X1 \o_values_reg[75][10]  (.D(o_values[10]), .CK(n_0_92), .Q(
      \o_values[75] [10]), .QN());
   DFF_X1 \o_values_reg[75][9]  (.D(o_values[9]), .CK(n_0_92), .Q(
      \o_values[75] [9]), .QN());
   DFF_X1 \o_values_reg[75][8]  (.D(o_values[8]), .CK(n_0_92), .Q(
      \o_values[75] [8]), .QN());
   DFF_X1 \o_values_reg[75][7]  (.D(o_values[7]), .CK(n_0_92), .Q(
      \o_values[75] [7]), .QN());
   DFF_X1 \o_values_reg[75][6]  (.D(o_values[6]), .CK(n_0_92), .Q(
      \o_values[75] [6]), .QN());
   DFF_X1 \o_values_reg[75][5]  (.D(o_values[5]), .CK(n_0_92), .Q(
      \o_values[75] [5]), .QN());
   DFF_X1 \o_values_reg[75][4]  (.D(o_values[4]), .CK(n_0_92), .Q(
      \o_values[75] [4]), .QN());
   DFF_X1 \o_values_reg[75][3]  (.D(o_values[3]), .CK(n_0_92), .Q(
      \o_values[75] [3]), .QN());
   DFF_X1 \o_values_reg[75][2]  (.D(o_values[2]), .CK(n_0_92), .Q(
      \o_values[75] [2]), .QN());
   DFF_X1 \o_values_reg[75][1]  (.D(o_values[1]), .CK(n_0_92), .Q(
      \o_values[75] [1]), .QN());
   DFF_X1 \o_values_reg[75][0]  (.D(o_values[0]), .CK(n_0_92), .Q(
      \o_values[75] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[74]_reg  (.CK(clk), .E(n_0_9), .SE(1'b0), 
      .GCK(n_0_93));
   DFF_X1 \o_values_reg[74][15]  (.D(o_values[15]), .CK(n_0_93), .Q(
      \o_values[74] [15]), .QN());
   DFF_X1 \o_values_reg[74][14]  (.D(o_values[14]), .CK(n_0_93), .Q(
      \o_values[74] [14]), .QN());
   DFF_X1 \o_values_reg[74][13]  (.D(o_values[13]), .CK(n_0_93), .Q(
      \o_values[74] [13]), .QN());
   DFF_X1 \o_values_reg[74][12]  (.D(o_values[12]), .CK(n_0_93), .Q(
      \o_values[74] [12]), .QN());
   DFF_X1 \o_values_reg[74][11]  (.D(o_values[11]), .CK(n_0_93), .Q(
      \o_values[74] [11]), .QN());
   DFF_X1 \o_values_reg[74][10]  (.D(o_values[10]), .CK(n_0_93), .Q(
      \o_values[74] [10]), .QN());
   DFF_X1 \o_values_reg[74][9]  (.D(o_values[9]), .CK(n_0_93), .Q(
      \o_values[74] [9]), .QN());
   DFF_X1 \o_values_reg[74][8]  (.D(o_values[8]), .CK(n_0_93), .Q(
      \o_values[74] [8]), .QN());
   DFF_X1 \o_values_reg[74][7]  (.D(o_values[7]), .CK(n_0_93), .Q(
      \o_values[74] [7]), .QN());
   DFF_X1 \o_values_reg[74][6]  (.D(o_values[6]), .CK(n_0_93), .Q(
      \o_values[74] [6]), .QN());
   DFF_X1 \o_values_reg[74][5]  (.D(o_values[5]), .CK(n_0_93), .Q(
      \o_values[74] [5]), .QN());
   DFF_X1 \o_values_reg[74][4]  (.D(o_values[4]), .CK(n_0_93), .Q(
      \o_values[74] [4]), .QN());
   DFF_X1 \o_values_reg[74][3]  (.D(o_values[3]), .CK(n_0_93), .Q(
      \o_values[74] [3]), .QN());
   DFF_X1 \o_values_reg[74][2]  (.D(o_values[2]), .CK(n_0_93), .Q(
      \o_values[74] [2]), .QN());
   DFF_X1 \o_values_reg[74][1]  (.D(o_values[1]), .CK(n_0_93), .Q(
      \o_values[74] [1]), .QN());
   DFF_X1 \o_values_reg[74][0]  (.D(o_values[0]), .CK(n_0_93), .Q(
      \o_values[74] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[73]_reg  (.CK(clk), .E(n_0_10), .SE(1'b0), 
      .GCK(n_0_94));
   DFF_X1 \o_values_reg[73][15]  (.D(o_values[15]), .CK(n_0_94), .Q(
      \o_values[73] [15]), .QN());
   DFF_X1 \o_values_reg[73][14]  (.D(o_values[14]), .CK(n_0_94), .Q(
      \o_values[73] [14]), .QN());
   DFF_X1 \o_values_reg[73][13]  (.D(o_values[13]), .CK(n_0_94), .Q(
      \o_values[73] [13]), .QN());
   DFF_X1 \o_values_reg[73][12]  (.D(o_values[12]), .CK(n_0_94), .Q(
      \o_values[73] [12]), .QN());
   DFF_X1 \o_values_reg[73][11]  (.D(o_values[11]), .CK(n_0_94), .Q(
      \o_values[73] [11]), .QN());
   DFF_X1 \o_values_reg[73][10]  (.D(o_values[10]), .CK(n_0_94), .Q(
      \o_values[73] [10]), .QN());
   DFF_X1 \o_values_reg[73][9]  (.D(o_values[9]), .CK(n_0_94), .Q(
      \o_values[73] [9]), .QN());
   DFF_X1 \o_values_reg[73][8]  (.D(o_values[8]), .CK(n_0_94), .Q(
      \o_values[73] [8]), .QN());
   DFF_X1 \o_values_reg[73][7]  (.D(o_values[7]), .CK(n_0_94), .Q(
      \o_values[73] [7]), .QN());
   DFF_X1 \o_values_reg[73][6]  (.D(o_values[6]), .CK(n_0_94), .Q(
      \o_values[73] [6]), .QN());
   DFF_X1 \o_values_reg[73][5]  (.D(o_values[5]), .CK(n_0_94), .Q(
      \o_values[73] [5]), .QN());
   DFF_X1 \o_values_reg[73][4]  (.D(o_values[4]), .CK(n_0_94), .Q(
      \o_values[73] [4]), .QN());
   DFF_X1 \o_values_reg[73][3]  (.D(o_values[3]), .CK(n_0_94), .Q(
      \o_values[73] [3]), .QN());
   DFF_X1 \o_values_reg[73][2]  (.D(o_values[2]), .CK(n_0_94), .Q(
      \o_values[73] [2]), .QN());
   DFF_X1 \o_values_reg[73][1]  (.D(o_values[1]), .CK(n_0_94), .Q(
      \o_values[73] [1]), .QN());
   DFF_X1 \o_values_reg[73][0]  (.D(o_values[0]), .CK(n_0_94), .Q(
      \o_values[73] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[72]_reg  (.CK(clk), .E(n_0_11), .SE(1'b0), 
      .GCK(n_0_95));
   DFF_X1 \o_values_reg[72][15]  (.D(o_values[15]), .CK(n_0_95), .Q(
      \o_values[72] [15]), .QN());
   DFF_X1 \o_values_reg[72][14]  (.D(o_values[14]), .CK(n_0_95), .Q(
      \o_values[72] [14]), .QN());
   DFF_X1 \o_values_reg[72][13]  (.D(o_values[13]), .CK(n_0_95), .Q(
      \o_values[72] [13]), .QN());
   DFF_X1 \o_values_reg[72][12]  (.D(o_values[12]), .CK(n_0_95), .Q(
      \o_values[72] [12]), .QN());
   DFF_X1 \o_values_reg[72][11]  (.D(o_values[11]), .CK(n_0_95), .Q(
      \o_values[72] [11]), .QN());
   DFF_X1 \o_values_reg[72][10]  (.D(o_values[10]), .CK(n_0_95), .Q(
      \o_values[72] [10]), .QN());
   DFF_X1 \o_values_reg[72][9]  (.D(o_values[9]), .CK(n_0_95), .Q(
      \o_values[72] [9]), .QN());
   DFF_X1 \o_values_reg[72][8]  (.D(o_values[8]), .CK(n_0_95), .Q(
      \o_values[72] [8]), .QN());
   DFF_X1 \o_values_reg[72][7]  (.D(o_values[7]), .CK(n_0_95), .Q(
      \o_values[72] [7]), .QN());
   DFF_X1 \o_values_reg[72][6]  (.D(o_values[6]), .CK(n_0_95), .Q(
      \o_values[72] [6]), .QN());
   DFF_X1 \o_values_reg[72][5]  (.D(o_values[5]), .CK(n_0_95), .Q(
      \o_values[72] [5]), .QN());
   DFF_X1 \o_values_reg[72][4]  (.D(o_values[4]), .CK(n_0_95), .Q(
      \o_values[72] [4]), .QN());
   DFF_X1 \o_values_reg[72][3]  (.D(o_values[3]), .CK(n_0_95), .Q(
      \o_values[72] [3]), .QN());
   DFF_X1 \o_values_reg[72][2]  (.D(o_values[2]), .CK(n_0_95), .Q(
      \o_values[72] [2]), .QN());
   DFF_X1 \o_values_reg[72][1]  (.D(o_values[1]), .CK(n_0_95), .Q(
      \o_values[72] [1]), .QN());
   DFF_X1 \o_values_reg[72][0]  (.D(o_values[0]), .CK(n_0_95), .Q(
      \o_values[72] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[71]_reg  (.CK(clk), .E(n_0_12), .SE(1'b0), 
      .GCK(n_0_96));
   DFF_X1 \o_values_reg[71][15]  (.D(o_values[15]), .CK(n_0_96), .Q(
      \o_values[71] [15]), .QN());
   DFF_X1 \o_values_reg[71][14]  (.D(o_values[14]), .CK(n_0_96), .Q(
      \o_values[71] [14]), .QN());
   DFF_X1 \o_values_reg[71][13]  (.D(o_values[13]), .CK(n_0_96), .Q(
      \o_values[71] [13]), .QN());
   DFF_X1 \o_values_reg[71][12]  (.D(o_values[12]), .CK(n_0_96), .Q(
      \o_values[71] [12]), .QN());
   DFF_X1 \o_values_reg[71][11]  (.D(o_values[11]), .CK(n_0_96), .Q(
      \o_values[71] [11]), .QN());
   DFF_X1 \o_values_reg[71][10]  (.D(o_values[10]), .CK(n_0_96), .Q(
      \o_values[71] [10]), .QN());
   DFF_X1 \o_values_reg[71][9]  (.D(o_values[9]), .CK(n_0_96), .Q(
      \o_values[71] [9]), .QN());
   DFF_X1 \o_values_reg[71][8]  (.D(o_values[8]), .CK(n_0_96), .Q(
      \o_values[71] [8]), .QN());
   DFF_X1 \o_values_reg[71][7]  (.D(o_values[7]), .CK(n_0_96), .Q(
      \o_values[71] [7]), .QN());
   DFF_X1 \o_values_reg[71][6]  (.D(o_values[6]), .CK(n_0_96), .Q(
      \o_values[71] [6]), .QN());
   DFF_X1 \o_values_reg[71][5]  (.D(o_values[5]), .CK(n_0_96), .Q(
      \o_values[71] [5]), .QN());
   DFF_X1 \o_values_reg[71][4]  (.D(o_values[4]), .CK(n_0_96), .Q(
      \o_values[71] [4]), .QN());
   DFF_X1 \o_values_reg[71][3]  (.D(o_values[3]), .CK(n_0_96), .Q(
      \o_values[71] [3]), .QN());
   DFF_X1 \o_values_reg[71][2]  (.D(o_values[2]), .CK(n_0_96), .Q(
      \o_values[71] [2]), .QN());
   DFF_X1 \o_values_reg[71][1]  (.D(o_values[1]), .CK(n_0_96), .Q(
      \o_values[71] [1]), .QN());
   DFF_X1 \o_values_reg[71][0]  (.D(o_values[0]), .CK(n_0_96), .Q(
      \o_values[71] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[70]_reg  (.CK(clk), .E(n_0_13), .SE(1'b0), 
      .GCK(n_0_97));
   DFF_X1 \o_values_reg[70][15]  (.D(o_values[15]), .CK(n_0_97), .Q(
      \o_values[70] [15]), .QN());
   DFF_X1 \o_values_reg[70][14]  (.D(o_values[14]), .CK(n_0_97), .Q(
      \o_values[70] [14]), .QN());
   DFF_X1 \o_values_reg[70][13]  (.D(o_values[13]), .CK(n_0_97), .Q(
      \o_values[70] [13]), .QN());
   DFF_X1 \o_values_reg[70][12]  (.D(o_values[12]), .CK(n_0_97), .Q(
      \o_values[70] [12]), .QN());
   DFF_X1 \o_values_reg[70][11]  (.D(o_values[11]), .CK(n_0_97), .Q(
      \o_values[70] [11]), .QN());
   DFF_X1 \o_values_reg[70][10]  (.D(o_values[10]), .CK(n_0_97), .Q(
      \o_values[70] [10]), .QN());
   DFF_X1 \o_values_reg[70][9]  (.D(o_values[9]), .CK(n_0_97), .Q(
      \o_values[70] [9]), .QN());
   DFF_X1 \o_values_reg[70][8]  (.D(o_values[8]), .CK(n_0_97), .Q(
      \o_values[70] [8]), .QN());
   DFF_X1 \o_values_reg[70][7]  (.D(o_values[7]), .CK(n_0_97), .Q(
      \o_values[70] [7]), .QN());
   DFF_X1 \o_values_reg[70][6]  (.D(o_values[6]), .CK(n_0_97), .Q(
      \o_values[70] [6]), .QN());
   DFF_X1 \o_values_reg[70][5]  (.D(o_values[5]), .CK(n_0_97), .Q(
      \o_values[70] [5]), .QN());
   DFF_X1 \o_values_reg[70][4]  (.D(o_values[4]), .CK(n_0_97), .Q(
      \o_values[70] [4]), .QN());
   DFF_X1 \o_values_reg[70][3]  (.D(o_values[3]), .CK(n_0_97), .Q(
      \o_values[70] [3]), .QN());
   DFF_X1 \o_values_reg[70][2]  (.D(o_values[2]), .CK(n_0_97), .Q(
      \o_values[70] [2]), .QN());
   DFF_X1 \o_values_reg[70][1]  (.D(o_values[1]), .CK(n_0_97), .Q(
      \o_values[70] [1]), .QN());
   DFF_X1 \o_values_reg[70][0]  (.D(o_values[0]), .CK(n_0_97), .Q(
      \o_values[70] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[69]_reg  (.CK(clk), .E(n_0_14), .SE(1'b0), 
      .GCK(n_0_98));
   DFF_X1 \o_values_reg[69][15]  (.D(o_values[15]), .CK(n_0_98), .Q(
      \o_values[69] [15]), .QN());
   DFF_X1 \o_values_reg[69][14]  (.D(o_values[14]), .CK(n_0_98), .Q(
      \o_values[69] [14]), .QN());
   DFF_X1 \o_values_reg[69][13]  (.D(o_values[13]), .CK(n_0_98), .Q(
      \o_values[69] [13]), .QN());
   DFF_X1 \o_values_reg[69][12]  (.D(o_values[12]), .CK(n_0_98), .Q(
      \o_values[69] [12]), .QN());
   DFF_X1 \o_values_reg[69][11]  (.D(o_values[11]), .CK(n_0_98), .Q(
      \o_values[69] [11]), .QN());
   DFF_X1 \o_values_reg[69][10]  (.D(o_values[10]), .CK(n_0_98), .Q(
      \o_values[69] [10]), .QN());
   DFF_X1 \o_values_reg[69][9]  (.D(o_values[9]), .CK(n_0_98), .Q(
      \o_values[69] [9]), .QN());
   DFF_X1 \o_values_reg[69][8]  (.D(o_values[8]), .CK(n_0_98), .Q(
      \o_values[69] [8]), .QN());
   DFF_X1 \o_values_reg[69][7]  (.D(o_values[7]), .CK(n_0_98), .Q(
      \o_values[69] [7]), .QN());
   DFF_X1 \o_values_reg[69][6]  (.D(o_values[6]), .CK(n_0_98), .Q(
      \o_values[69] [6]), .QN());
   DFF_X1 \o_values_reg[69][5]  (.D(o_values[5]), .CK(n_0_98), .Q(
      \o_values[69] [5]), .QN());
   DFF_X1 \o_values_reg[69][4]  (.D(o_values[4]), .CK(n_0_98), .Q(
      \o_values[69] [4]), .QN());
   DFF_X1 \o_values_reg[69][3]  (.D(o_values[3]), .CK(n_0_98), .Q(
      \o_values[69] [3]), .QN());
   DFF_X1 \o_values_reg[69][2]  (.D(o_values[2]), .CK(n_0_98), .Q(
      \o_values[69] [2]), .QN());
   DFF_X1 \o_values_reg[69][1]  (.D(o_values[1]), .CK(n_0_98), .Q(
      \o_values[69] [1]), .QN());
   DFF_X1 \o_values_reg[69][0]  (.D(o_values[0]), .CK(n_0_98), .Q(
      \o_values[69] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[68]_reg  (.CK(clk), .E(n_0_15), .SE(1'b0), 
      .GCK(n_0_99));
   DFF_X1 \o_values_reg[68][15]  (.D(o_values[15]), .CK(n_0_99), .Q(
      \o_values[68] [15]), .QN());
   DFF_X1 \o_values_reg[68][14]  (.D(o_values[14]), .CK(n_0_99), .Q(
      \o_values[68] [14]), .QN());
   DFF_X1 \o_values_reg[68][13]  (.D(o_values[13]), .CK(n_0_99), .Q(
      \o_values[68] [13]), .QN());
   DFF_X1 \o_values_reg[68][12]  (.D(o_values[12]), .CK(n_0_99), .Q(
      \o_values[68] [12]), .QN());
   DFF_X1 \o_values_reg[68][11]  (.D(o_values[11]), .CK(n_0_99), .Q(
      \o_values[68] [11]), .QN());
   DFF_X1 \o_values_reg[68][10]  (.D(o_values[10]), .CK(n_0_99), .Q(
      \o_values[68] [10]), .QN());
   DFF_X1 \o_values_reg[68][9]  (.D(o_values[9]), .CK(n_0_99), .Q(
      \o_values[68] [9]), .QN());
   DFF_X1 \o_values_reg[68][8]  (.D(o_values[8]), .CK(n_0_99), .Q(
      \o_values[68] [8]), .QN());
   DFF_X1 \o_values_reg[68][7]  (.D(o_values[7]), .CK(n_0_99), .Q(
      \o_values[68] [7]), .QN());
   DFF_X1 \o_values_reg[68][6]  (.D(o_values[6]), .CK(n_0_99), .Q(
      \o_values[68] [6]), .QN());
   DFF_X1 \o_values_reg[68][5]  (.D(o_values[5]), .CK(n_0_99), .Q(
      \o_values[68] [5]), .QN());
   DFF_X1 \o_values_reg[68][4]  (.D(o_values[4]), .CK(n_0_99), .Q(
      \o_values[68] [4]), .QN());
   DFF_X1 \o_values_reg[68][3]  (.D(o_values[3]), .CK(n_0_99), .Q(
      \o_values[68] [3]), .QN());
   DFF_X1 \o_values_reg[68][2]  (.D(o_values[2]), .CK(n_0_99), .Q(
      \o_values[68] [2]), .QN());
   DFF_X1 \o_values_reg[68][1]  (.D(o_values[1]), .CK(n_0_99), .Q(
      \o_values[68] [1]), .QN());
   DFF_X1 \o_values_reg[68][0]  (.D(o_values[0]), .CK(n_0_99), .Q(
      \o_values[68] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[67]_reg  (.CK(clk), .E(n_0_16), .SE(1'b0), 
      .GCK(n_0_100));
   DFF_X1 \o_values_reg[67][15]  (.D(o_values[15]), .CK(n_0_100), .Q(
      \o_values[67] [15]), .QN());
   DFF_X1 \o_values_reg[67][14]  (.D(o_values[14]), .CK(n_0_100), .Q(
      \o_values[67] [14]), .QN());
   DFF_X1 \o_values_reg[67][13]  (.D(o_values[13]), .CK(n_0_100), .Q(
      \o_values[67] [13]), .QN());
   DFF_X1 \o_values_reg[67][12]  (.D(o_values[12]), .CK(n_0_100), .Q(
      \o_values[67] [12]), .QN());
   DFF_X1 \o_values_reg[67][11]  (.D(o_values[11]), .CK(n_0_100), .Q(
      \o_values[67] [11]), .QN());
   DFF_X1 \o_values_reg[67][10]  (.D(o_values[10]), .CK(n_0_100), .Q(
      \o_values[67] [10]), .QN());
   DFF_X1 \o_values_reg[67][9]  (.D(o_values[9]), .CK(n_0_100), .Q(
      \o_values[67] [9]), .QN());
   DFF_X1 \o_values_reg[67][8]  (.D(o_values[8]), .CK(n_0_100), .Q(
      \o_values[67] [8]), .QN());
   DFF_X1 \o_values_reg[67][7]  (.D(o_values[7]), .CK(n_0_100), .Q(
      \o_values[67] [7]), .QN());
   DFF_X1 \o_values_reg[67][6]  (.D(o_values[6]), .CK(n_0_100), .Q(
      \o_values[67] [6]), .QN());
   DFF_X1 \o_values_reg[67][5]  (.D(o_values[5]), .CK(n_0_100), .Q(
      \o_values[67] [5]), .QN());
   DFF_X1 \o_values_reg[67][4]  (.D(o_values[4]), .CK(n_0_100), .Q(
      \o_values[67] [4]), .QN());
   DFF_X1 \o_values_reg[67][3]  (.D(o_values[3]), .CK(n_0_100), .Q(
      \o_values[67] [3]), .QN());
   DFF_X1 \o_values_reg[67][2]  (.D(o_values[2]), .CK(n_0_100), .Q(
      \o_values[67] [2]), .QN());
   DFF_X1 \o_values_reg[67][1]  (.D(o_values[1]), .CK(n_0_100), .Q(
      \o_values[67] [1]), .QN());
   DFF_X1 \o_values_reg[67][0]  (.D(o_values[0]), .CK(n_0_100), .Q(
      \o_values[67] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[66]_reg  (.CK(clk), .E(n_0_17), .SE(1'b0), 
      .GCK(n_0_101));
   DFF_X1 \o_values_reg[66][15]  (.D(o_values[15]), .CK(n_0_101), .Q(
      \o_values[66] [15]), .QN());
   DFF_X1 \o_values_reg[66][14]  (.D(o_values[14]), .CK(n_0_101), .Q(
      \o_values[66] [14]), .QN());
   DFF_X1 \o_values_reg[66][13]  (.D(o_values[13]), .CK(n_0_101), .Q(
      \o_values[66] [13]), .QN());
   DFF_X1 \o_values_reg[66][12]  (.D(o_values[12]), .CK(n_0_101), .Q(
      \o_values[66] [12]), .QN());
   DFF_X1 \o_values_reg[66][11]  (.D(o_values[11]), .CK(n_0_101), .Q(
      \o_values[66] [11]), .QN());
   DFF_X1 \o_values_reg[66][10]  (.D(o_values[10]), .CK(n_0_101), .Q(
      \o_values[66] [10]), .QN());
   DFF_X1 \o_values_reg[66][9]  (.D(o_values[9]), .CK(n_0_101), .Q(
      \o_values[66] [9]), .QN());
   DFF_X1 \o_values_reg[66][8]  (.D(o_values[8]), .CK(n_0_101), .Q(
      \o_values[66] [8]), .QN());
   DFF_X1 \o_values_reg[66][7]  (.D(o_values[7]), .CK(n_0_101), .Q(
      \o_values[66] [7]), .QN());
   DFF_X1 \o_values_reg[66][6]  (.D(o_values[6]), .CK(n_0_101), .Q(
      \o_values[66] [6]), .QN());
   DFF_X1 \o_values_reg[66][5]  (.D(o_values[5]), .CK(n_0_101), .Q(
      \o_values[66] [5]), .QN());
   DFF_X1 \o_values_reg[66][4]  (.D(o_values[4]), .CK(n_0_101), .Q(
      \o_values[66] [4]), .QN());
   DFF_X1 \o_values_reg[66][3]  (.D(o_values[3]), .CK(n_0_101), .Q(
      \o_values[66] [3]), .QN());
   DFF_X1 \o_values_reg[66][2]  (.D(o_values[2]), .CK(n_0_101), .Q(
      \o_values[66] [2]), .QN());
   DFF_X1 \o_values_reg[66][1]  (.D(o_values[1]), .CK(n_0_101), .Q(
      \o_values[66] [1]), .QN());
   DFF_X1 \o_values_reg[66][0]  (.D(o_values[0]), .CK(n_0_101), .Q(
      \o_values[66] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[65]_reg  (.CK(clk), .E(n_0_18), .SE(1'b0), 
      .GCK(n_0_102));
   DFF_X1 \o_values_reg[65][15]  (.D(o_values[15]), .CK(n_0_102), .Q(
      \o_values[65] [15]), .QN());
   DFF_X1 \o_values_reg[65][14]  (.D(o_values[14]), .CK(n_0_102), .Q(
      \o_values[65] [14]), .QN());
   DFF_X1 \o_values_reg[65][13]  (.D(o_values[13]), .CK(n_0_102), .Q(
      \o_values[65] [13]), .QN());
   DFF_X1 \o_values_reg[65][12]  (.D(o_values[12]), .CK(n_0_102), .Q(
      \o_values[65] [12]), .QN());
   DFF_X1 \o_values_reg[65][11]  (.D(o_values[11]), .CK(n_0_102), .Q(
      \o_values[65] [11]), .QN());
   DFF_X1 \o_values_reg[65][10]  (.D(o_values[10]), .CK(n_0_102), .Q(
      \o_values[65] [10]), .QN());
   DFF_X1 \o_values_reg[65][9]  (.D(o_values[9]), .CK(n_0_102), .Q(
      \o_values[65] [9]), .QN());
   DFF_X1 \o_values_reg[65][8]  (.D(o_values[8]), .CK(n_0_102), .Q(
      \o_values[65] [8]), .QN());
   DFF_X1 \o_values_reg[65][7]  (.D(o_values[7]), .CK(n_0_102), .Q(
      \o_values[65] [7]), .QN());
   DFF_X1 \o_values_reg[65][6]  (.D(o_values[6]), .CK(n_0_102), .Q(
      \o_values[65] [6]), .QN());
   DFF_X1 \o_values_reg[65][5]  (.D(o_values[5]), .CK(n_0_102), .Q(
      \o_values[65] [5]), .QN());
   DFF_X1 \o_values_reg[65][4]  (.D(o_values[4]), .CK(n_0_102), .Q(
      \o_values[65] [4]), .QN());
   DFF_X1 \o_values_reg[65][3]  (.D(o_values[3]), .CK(n_0_102), .Q(
      \o_values[65] [3]), .QN());
   DFF_X1 \o_values_reg[65][2]  (.D(o_values[2]), .CK(n_0_102), .Q(
      \o_values[65] [2]), .QN());
   DFF_X1 \o_values_reg[65][1]  (.D(o_values[1]), .CK(n_0_102), .Q(
      \o_values[65] [1]), .QN());
   DFF_X1 \o_values_reg[65][0]  (.D(o_values[0]), .CK(n_0_102), .Q(
      \o_values[65] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[64]_reg  (.CK(clk), .E(n_0_19), .SE(1'b0), 
      .GCK(n_0_103));
   DFF_X1 \o_values_reg[64][15]  (.D(o_values[15]), .CK(n_0_103), .Q(
      \o_values[64] [15]), .QN());
   DFF_X1 \o_values_reg[64][14]  (.D(o_values[14]), .CK(n_0_103), .Q(
      \o_values[64] [14]), .QN());
   DFF_X1 \o_values_reg[64][13]  (.D(o_values[13]), .CK(n_0_103), .Q(
      \o_values[64] [13]), .QN());
   DFF_X1 \o_values_reg[64][12]  (.D(o_values[12]), .CK(n_0_103), .Q(
      \o_values[64] [12]), .QN());
   DFF_X1 \o_values_reg[64][11]  (.D(o_values[11]), .CK(n_0_103), .Q(
      \o_values[64] [11]), .QN());
   DFF_X1 \o_values_reg[64][10]  (.D(o_values[10]), .CK(n_0_103), .Q(
      \o_values[64] [10]), .QN());
   DFF_X1 \o_values_reg[64][9]  (.D(o_values[9]), .CK(n_0_103), .Q(
      \o_values[64] [9]), .QN());
   DFF_X1 \o_values_reg[64][8]  (.D(o_values[8]), .CK(n_0_103), .Q(
      \o_values[64] [8]), .QN());
   DFF_X1 \o_values_reg[64][7]  (.D(o_values[7]), .CK(n_0_103), .Q(
      \o_values[64] [7]), .QN());
   DFF_X1 \o_values_reg[64][6]  (.D(o_values[6]), .CK(n_0_103), .Q(
      \o_values[64] [6]), .QN());
   DFF_X1 \o_values_reg[64][5]  (.D(o_values[5]), .CK(n_0_103), .Q(
      \o_values[64] [5]), .QN());
   DFF_X1 \o_values_reg[64][4]  (.D(o_values[4]), .CK(n_0_103), .Q(
      \o_values[64] [4]), .QN());
   DFF_X1 \o_values_reg[64][3]  (.D(o_values[3]), .CK(n_0_103), .Q(
      \o_values[64] [3]), .QN());
   DFF_X1 \o_values_reg[64][2]  (.D(o_values[2]), .CK(n_0_103), .Q(
      \o_values[64] [2]), .QN());
   DFF_X1 \o_values_reg[64][1]  (.D(o_values[1]), .CK(n_0_103), .Q(
      \o_values[64] [1]), .QN());
   DFF_X1 \o_values_reg[64][0]  (.D(o_values[0]), .CK(n_0_103), .Q(
      \o_values[64] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[63]_reg  (.CK(clk), .E(n_0_20), .SE(1'b0), 
      .GCK(n_0_104));
   DFF_X1 \o_values_reg[63][15]  (.D(o_values[15]), .CK(n_0_104), .Q(
      \o_values[63] [15]), .QN());
   DFF_X1 \o_values_reg[63][14]  (.D(o_values[14]), .CK(n_0_104), .Q(
      \o_values[63] [14]), .QN());
   DFF_X1 \o_values_reg[63][13]  (.D(o_values[13]), .CK(n_0_104), .Q(
      \o_values[63] [13]), .QN());
   DFF_X1 \o_values_reg[63][12]  (.D(o_values[12]), .CK(n_0_104), .Q(
      \o_values[63] [12]), .QN());
   DFF_X1 \o_values_reg[63][11]  (.D(o_values[11]), .CK(n_0_104), .Q(
      \o_values[63] [11]), .QN());
   DFF_X1 \o_values_reg[63][10]  (.D(o_values[10]), .CK(n_0_104), .Q(
      \o_values[63] [10]), .QN());
   DFF_X1 \o_values_reg[63][9]  (.D(o_values[9]), .CK(n_0_104), .Q(
      \o_values[63] [9]), .QN());
   DFF_X1 \o_values_reg[63][8]  (.D(o_values[8]), .CK(n_0_104), .Q(
      \o_values[63] [8]), .QN());
   DFF_X1 \o_values_reg[63][7]  (.D(o_values[7]), .CK(n_0_104), .Q(
      \o_values[63] [7]), .QN());
   DFF_X1 \o_values_reg[63][6]  (.D(o_values[6]), .CK(n_0_104), .Q(
      \o_values[63] [6]), .QN());
   DFF_X1 \o_values_reg[63][5]  (.D(o_values[5]), .CK(n_0_104), .Q(
      \o_values[63] [5]), .QN());
   DFF_X1 \o_values_reg[63][4]  (.D(o_values[4]), .CK(n_0_104), .Q(
      \o_values[63] [4]), .QN());
   DFF_X1 \o_values_reg[63][3]  (.D(o_values[3]), .CK(n_0_104), .Q(
      \o_values[63] [3]), .QN());
   DFF_X1 \o_values_reg[63][2]  (.D(o_values[2]), .CK(n_0_104), .Q(
      \o_values[63] [2]), .QN());
   DFF_X1 \o_values_reg[63][1]  (.D(o_values[1]), .CK(n_0_104), .Q(
      \o_values[63] [1]), .QN());
   DFF_X1 \o_values_reg[63][0]  (.D(o_values[0]), .CK(n_0_104), .Q(
      \o_values[63] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[62]_reg  (.CK(clk), .E(n_0_21), .SE(1'b0), 
      .GCK(n_0_105));
   DFF_X1 \o_values_reg[62][15]  (.D(o_values[15]), .CK(n_0_105), .Q(
      \o_values[62] [15]), .QN());
   DFF_X1 \o_values_reg[62][14]  (.D(o_values[14]), .CK(n_0_105), .Q(
      \o_values[62] [14]), .QN());
   DFF_X1 \o_values_reg[62][13]  (.D(o_values[13]), .CK(n_0_105), .Q(
      \o_values[62] [13]), .QN());
   DFF_X1 \o_values_reg[62][12]  (.D(o_values[12]), .CK(n_0_105), .Q(
      \o_values[62] [12]), .QN());
   DFF_X1 \o_values_reg[62][11]  (.D(o_values[11]), .CK(n_0_105), .Q(
      \o_values[62] [11]), .QN());
   DFF_X1 \o_values_reg[62][10]  (.D(o_values[10]), .CK(n_0_105), .Q(
      \o_values[62] [10]), .QN());
   DFF_X1 \o_values_reg[62][9]  (.D(o_values[9]), .CK(n_0_105), .Q(
      \o_values[62] [9]), .QN());
   DFF_X1 \o_values_reg[62][8]  (.D(o_values[8]), .CK(n_0_105), .Q(
      \o_values[62] [8]), .QN());
   DFF_X1 \o_values_reg[62][7]  (.D(o_values[7]), .CK(n_0_105), .Q(
      \o_values[62] [7]), .QN());
   DFF_X1 \o_values_reg[62][6]  (.D(o_values[6]), .CK(n_0_105), .Q(
      \o_values[62] [6]), .QN());
   DFF_X1 \o_values_reg[62][5]  (.D(o_values[5]), .CK(n_0_105), .Q(
      \o_values[62] [5]), .QN());
   DFF_X1 \o_values_reg[62][4]  (.D(o_values[4]), .CK(n_0_105), .Q(
      \o_values[62] [4]), .QN());
   DFF_X1 \o_values_reg[62][3]  (.D(o_values[3]), .CK(n_0_105), .Q(
      \o_values[62] [3]), .QN());
   DFF_X1 \o_values_reg[62][2]  (.D(o_values[2]), .CK(n_0_105), .Q(
      \o_values[62] [2]), .QN());
   DFF_X1 \o_values_reg[62][1]  (.D(o_values[1]), .CK(n_0_105), .Q(
      \o_values[62] [1]), .QN());
   DFF_X1 \o_values_reg[62][0]  (.D(o_values[0]), .CK(n_0_105), .Q(
      \o_values[62] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[61]_reg  (.CK(clk), .E(n_0_22), .SE(1'b0), 
      .GCK(n_0_106));
   DFF_X1 \o_values_reg[61][15]  (.D(o_values[15]), .CK(n_0_106), .Q(
      \o_values[61] [15]), .QN());
   DFF_X1 \o_values_reg[61][14]  (.D(o_values[14]), .CK(n_0_106), .Q(
      \o_values[61] [14]), .QN());
   DFF_X1 \o_values_reg[61][13]  (.D(o_values[13]), .CK(n_0_106), .Q(
      \o_values[61] [13]), .QN());
   DFF_X1 \o_values_reg[61][12]  (.D(o_values[12]), .CK(n_0_106), .Q(
      \o_values[61] [12]), .QN());
   DFF_X1 \o_values_reg[61][11]  (.D(o_values[11]), .CK(n_0_106), .Q(
      \o_values[61] [11]), .QN());
   DFF_X1 \o_values_reg[61][10]  (.D(o_values[10]), .CK(n_0_106), .Q(
      \o_values[61] [10]), .QN());
   DFF_X1 \o_values_reg[61][9]  (.D(o_values[9]), .CK(n_0_106), .Q(
      \o_values[61] [9]), .QN());
   DFF_X1 \o_values_reg[61][8]  (.D(o_values[8]), .CK(n_0_106), .Q(
      \o_values[61] [8]), .QN());
   DFF_X1 \o_values_reg[61][7]  (.D(o_values[7]), .CK(n_0_106), .Q(
      \o_values[61] [7]), .QN());
   DFF_X1 \o_values_reg[61][6]  (.D(o_values[6]), .CK(n_0_106), .Q(
      \o_values[61] [6]), .QN());
   DFF_X1 \o_values_reg[61][5]  (.D(o_values[5]), .CK(n_0_106), .Q(
      \o_values[61] [5]), .QN());
   DFF_X1 \o_values_reg[61][4]  (.D(o_values[4]), .CK(n_0_106), .Q(
      \o_values[61] [4]), .QN());
   DFF_X1 \o_values_reg[61][3]  (.D(o_values[3]), .CK(n_0_106), .Q(
      \o_values[61] [3]), .QN());
   DFF_X1 \o_values_reg[61][2]  (.D(o_values[2]), .CK(n_0_106), .Q(
      \o_values[61] [2]), .QN());
   DFF_X1 \o_values_reg[61][1]  (.D(o_values[1]), .CK(n_0_106), .Q(
      \o_values[61] [1]), .QN());
   DFF_X1 \o_values_reg[61][0]  (.D(o_values[0]), .CK(n_0_106), .Q(
      \o_values[61] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[60]_reg  (.CK(clk), .E(n_0_23), .SE(1'b0), 
      .GCK(n_0_107));
   DFF_X1 \o_values_reg[60][15]  (.D(o_values[15]), .CK(n_0_107), .Q(
      \o_values[60] [15]), .QN());
   DFF_X1 \o_values_reg[60][14]  (.D(o_values[14]), .CK(n_0_107), .Q(
      \o_values[60] [14]), .QN());
   DFF_X1 \o_values_reg[60][13]  (.D(o_values[13]), .CK(n_0_107), .Q(
      \o_values[60] [13]), .QN());
   DFF_X1 \o_values_reg[60][12]  (.D(o_values[12]), .CK(n_0_107), .Q(
      \o_values[60] [12]), .QN());
   DFF_X1 \o_values_reg[60][11]  (.D(o_values[11]), .CK(n_0_107), .Q(
      \o_values[60] [11]), .QN());
   DFF_X1 \o_values_reg[60][10]  (.D(o_values[10]), .CK(n_0_107), .Q(
      \o_values[60] [10]), .QN());
   DFF_X1 \o_values_reg[60][9]  (.D(o_values[9]), .CK(n_0_107), .Q(
      \o_values[60] [9]), .QN());
   DFF_X1 \o_values_reg[60][8]  (.D(o_values[8]), .CK(n_0_107), .Q(
      \o_values[60] [8]), .QN());
   DFF_X1 \o_values_reg[60][7]  (.D(o_values[7]), .CK(n_0_107), .Q(
      \o_values[60] [7]), .QN());
   DFF_X1 \o_values_reg[60][6]  (.D(o_values[6]), .CK(n_0_107), .Q(
      \o_values[60] [6]), .QN());
   DFF_X1 \o_values_reg[60][5]  (.D(o_values[5]), .CK(n_0_107), .Q(
      \o_values[60] [5]), .QN());
   DFF_X1 \o_values_reg[60][4]  (.D(o_values[4]), .CK(n_0_107), .Q(
      \o_values[60] [4]), .QN());
   DFF_X1 \o_values_reg[60][3]  (.D(o_values[3]), .CK(n_0_107), .Q(
      \o_values[60] [3]), .QN());
   DFF_X1 \o_values_reg[60][2]  (.D(o_values[2]), .CK(n_0_107), .Q(
      \o_values[60] [2]), .QN());
   DFF_X1 \o_values_reg[60][1]  (.D(o_values[1]), .CK(n_0_107), .Q(
      \o_values[60] [1]), .QN());
   DFF_X1 \o_values_reg[60][0]  (.D(o_values[0]), .CK(n_0_107), .Q(
      \o_values[60] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[59]_reg  (.CK(clk), .E(n_0_24), .SE(1'b0), 
      .GCK(n_0_108));
   DFF_X1 \o_values_reg[59][15]  (.D(o_values[15]), .CK(n_0_108), .Q(
      \o_values[59] [15]), .QN());
   DFF_X1 \o_values_reg[59][14]  (.D(o_values[14]), .CK(n_0_108), .Q(
      \o_values[59] [14]), .QN());
   DFF_X1 \o_values_reg[59][13]  (.D(o_values[13]), .CK(n_0_108), .Q(
      \o_values[59] [13]), .QN());
   DFF_X1 \o_values_reg[59][12]  (.D(o_values[12]), .CK(n_0_108), .Q(
      \o_values[59] [12]), .QN());
   DFF_X1 \o_values_reg[59][11]  (.D(o_values[11]), .CK(n_0_108), .Q(
      \o_values[59] [11]), .QN());
   DFF_X1 \o_values_reg[59][10]  (.D(o_values[10]), .CK(n_0_108), .Q(
      \o_values[59] [10]), .QN());
   DFF_X1 \o_values_reg[59][9]  (.D(o_values[9]), .CK(n_0_108), .Q(
      \o_values[59] [9]), .QN());
   DFF_X1 \o_values_reg[59][8]  (.D(o_values[8]), .CK(n_0_108), .Q(
      \o_values[59] [8]), .QN());
   DFF_X1 \o_values_reg[59][7]  (.D(o_values[7]), .CK(n_0_108), .Q(
      \o_values[59] [7]), .QN());
   DFF_X1 \o_values_reg[59][6]  (.D(o_values[6]), .CK(n_0_108), .Q(
      \o_values[59] [6]), .QN());
   DFF_X1 \o_values_reg[59][5]  (.D(o_values[5]), .CK(n_0_108), .Q(
      \o_values[59] [5]), .QN());
   DFF_X1 \o_values_reg[59][4]  (.D(o_values[4]), .CK(n_0_108), .Q(
      \o_values[59] [4]), .QN());
   DFF_X1 \o_values_reg[59][3]  (.D(o_values[3]), .CK(n_0_108), .Q(
      \o_values[59] [3]), .QN());
   DFF_X1 \o_values_reg[59][2]  (.D(o_values[2]), .CK(n_0_108), .Q(
      \o_values[59] [2]), .QN());
   DFF_X1 \o_values_reg[59][1]  (.D(o_values[1]), .CK(n_0_108), .Q(
      \o_values[59] [1]), .QN());
   DFF_X1 \o_values_reg[59][0]  (.D(o_values[0]), .CK(n_0_108), .Q(
      \o_values[59] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[58]_reg  (.CK(clk), .E(n_0_25), .SE(1'b0), 
      .GCK(n_0_109));
   DFF_X1 \o_values_reg[58][15]  (.D(o_values[15]), .CK(n_0_109), .Q(
      \o_values[58] [15]), .QN());
   DFF_X1 \o_values_reg[58][14]  (.D(o_values[14]), .CK(n_0_109), .Q(
      \o_values[58] [14]), .QN());
   DFF_X1 \o_values_reg[58][13]  (.D(o_values[13]), .CK(n_0_109), .Q(
      \o_values[58] [13]), .QN());
   DFF_X1 \o_values_reg[58][12]  (.D(o_values[12]), .CK(n_0_109), .Q(
      \o_values[58] [12]), .QN());
   DFF_X1 \o_values_reg[58][11]  (.D(o_values[11]), .CK(n_0_109), .Q(
      \o_values[58] [11]), .QN());
   DFF_X1 \o_values_reg[58][10]  (.D(o_values[10]), .CK(n_0_109), .Q(
      \o_values[58] [10]), .QN());
   DFF_X1 \o_values_reg[58][9]  (.D(o_values[9]), .CK(n_0_109), .Q(
      \o_values[58] [9]), .QN());
   DFF_X1 \o_values_reg[58][8]  (.D(o_values[8]), .CK(n_0_109), .Q(
      \o_values[58] [8]), .QN());
   DFF_X1 \o_values_reg[58][7]  (.D(o_values[7]), .CK(n_0_109), .Q(
      \o_values[58] [7]), .QN());
   DFF_X1 \o_values_reg[58][6]  (.D(o_values[6]), .CK(n_0_109), .Q(
      \o_values[58] [6]), .QN());
   DFF_X1 \o_values_reg[58][5]  (.D(o_values[5]), .CK(n_0_109), .Q(
      \o_values[58] [5]), .QN());
   DFF_X1 \o_values_reg[58][4]  (.D(o_values[4]), .CK(n_0_109), .Q(
      \o_values[58] [4]), .QN());
   DFF_X1 \o_values_reg[58][3]  (.D(o_values[3]), .CK(n_0_109), .Q(
      \o_values[58] [3]), .QN());
   DFF_X1 \o_values_reg[58][2]  (.D(o_values[2]), .CK(n_0_109), .Q(
      \o_values[58] [2]), .QN());
   DFF_X1 \o_values_reg[58][1]  (.D(o_values[1]), .CK(n_0_109), .Q(
      \o_values[58] [1]), .QN());
   DFF_X1 \o_values_reg[58][0]  (.D(o_values[0]), .CK(n_0_109), .Q(
      \o_values[58] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[57]_reg  (.CK(clk), .E(n_0_26), .SE(1'b0), 
      .GCK(n_0_110));
   DFF_X1 \o_values_reg[57][15]  (.D(o_values[15]), .CK(n_0_110), .Q(
      \o_values[57] [15]), .QN());
   DFF_X1 \o_values_reg[57][14]  (.D(o_values[14]), .CK(n_0_110), .Q(
      \o_values[57] [14]), .QN());
   DFF_X1 \o_values_reg[57][13]  (.D(o_values[13]), .CK(n_0_110), .Q(
      \o_values[57] [13]), .QN());
   DFF_X1 \o_values_reg[57][12]  (.D(o_values[12]), .CK(n_0_110), .Q(
      \o_values[57] [12]), .QN());
   DFF_X1 \o_values_reg[57][11]  (.D(o_values[11]), .CK(n_0_110), .Q(
      \o_values[57] [11]), .QN());
   DFF_X1 \o_values_reg[57][10]  (.D(o_values[10]), .CK(n_0_110), .Q(
      \o_values[57] [10]), .QN());
   DFF_X1 \o_values_reg[57][9]  (.D(o_values[9]), .CK(n_0_110), .Q(
      \o_values[57] [9]), .QN());
   DFF_X1 \o_values_reg[57][8]  (.D(o_values[8]), .CK(n_0_110), .Q(
      \o_values[57] [8]), .QN());
   DFF_X1 \o_values_reg[57][7]  (.D(o_values[7]), .CK(n_0_110), .Q(
      \o_values[57] [7]), .QN());
   DFF_X1 \o_values_reg[57][6]  (.D(o_values[6]), .CK(n_0_110), .Q(
      \o_values[57] [6]), .QN());
   DFF_X1 \o_values_reg[57][5]  (.D(o_values[5]), .CK(n_0_110), .Q(
      \o_values[57] [5]), .QN());
   DFF_X1 \o_values_reg[57][4]  (.D(o_values[4]), .CK(n_0_110), .Q(
      \o_values[57] [4]), .QN());
   DFF_X1 \o_values_reg[57][3]  (.D(o_values[3]), .CK(n_0_110), .Q(
      \o_values[57] [3]), .QN());
   DFF_X1 \o_values_reg[57][2]  (.D(o_values[2]), .CK(n_0_110), .Q(
      \o_values[57] [2]), .QN());
   DFF_X1 \o_values_reg[57][1]  (.D(o_values[1]), .CK(n_0_110), .Q(
      \o_values[57] [1]), .QN());
   DFF_X1 \o_values_reg[57][0]  (.D(o_values[0]), .CK(n_0_110), .Q(
      \o_values[57] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[56]_reg  (.CK(clk), .E(n_0_27), .SE(1'b0), 
      .GCK(n_0_111));
   DFF_X1 \o_values_reg[56][15]  (.D(o_values[15]), .CK(n_0_111), .Q(
      \o_values[56] [15]), .QN());
   DFF_X1 \o_values_reg[56][14]  (.D(o_values[14]), .CK(n_0_111), .Q(
      \o_values[56] [14]), .QN());
   DFF_X1 \o_values_reg[56][13]  (.D(o_values[13]), .CK(n_0_111), .Q(
      \o_values[56] [13]), .QN());
   DFF_X1 \o_values_reg[56][12]  (.D(o_values[12]), .CK(n_0_111), .Q(
      \o_values[56] [12]), .QN());
   DFF_X1 \o_values_reg[56][11]  (.D(o_values[11]), .CK(n_0_111), .Q(
      \o_values[56] [11]), .QN());
   DFF_X1 \o_values_reg[56][10]  (.D(o_values[10]), .CK(n_0_111), .Q(
      \o_values[56] [10]), .QN());
   DFF_X1 \o_values_reg[56][9]  (.D(o_values[9]), .CK(n_0_111), .Q(
      \o_values[56] [9]), .QN());
   DFF_X1 \o_values_reg[56][8]  (.D(o_values[8]), .CK(n_0_111), .Q(
      \o_values[56] [8]), .QN());
   DFF_X1 \o_values_reg[56][7]  (.D(o_values[7]), .CK(n_0_111), .Q(
      \o_values[56] [7]), .QN());
   DFF_X1 \o_values_reg[56][6]  (.D(o_values[6]), .CK(n_0_111), .Q(
      \o_values[56] [6]), .QN());
   DFF_X1 \o_values_reg[56][5]  (.D(o_values[5]), .CK(n_0_111), .Q(
      \o_values[56] [5]), .QN());
   DFF_X1 \o_values_reg[56][4]  (.D(o_values[4]), .CK(n_0_111), .Q(
      \o_values[56] [4]), .QN());
   DFF_X1 \o_values_reg[56][3]  (.D(o_values[3]), .CK(n_0_111), .Q(
      \o_values[56] [3]), .QN());
   DFF_X1 \o_values_reg[56][2]  (.D(o_values[2]), .CK(n_0_111), .Q(
      \o_values[56] [2]), .QN());
   DFF_X1 \o_values_reg[56][1]  (.D(o_values[1]), .CK(n_0_111), .Q(
      \o_values[56] [1]), .QN());
   DFF_X1 \o_values_reg[56][0]  (.D(o_values[0]), .CK(n_0_111), .Q(
      \o_values[56] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[55]_reg  (.CK(clk), .E(n_0_28), .SE(1'b0), 
      .GCK(n_0_112));
   DFF_X1 \o_values_reg[55][15]  (.D(o_values[15]), .CK(n_0_112), .Q(
      \o_values[55] [15]), .QN());
   DFF_X1 \o_values_reg[55][14]  (.D(o_values[14]), .CK(n_0_112), .Q(
      \o_values[55] [14]), .QN());
   DFF_X1 \o_values_reg[55][13]  (.D(o_values[13]), .CK(n_0_112), .Q(
      \o_values[55] [13]), .QN());
   DFF_X1 \o_values_reg[55][12]  (.D(o_values[12]), .CK(n_0_112), .Q(
      \o_values[55] [12]), .QN());
   DFF_X1 \o_values_reg[55][11]  (.D(o_values[11]), .CK(n_0_112), .Q(
      \o_values[55] [11]), .QN());
   DFF_X1 \o_values_reg[55][10]  (.D(o_values[10]), .CK(n_0_112), .Q(
      \o_values[55] [10]), .QN());
   DFF_X1 \o_values_reg[55][9]  (.D(o_values[9]), .CK(n_0_112), .Q(
      \o_values[55] [9]), .QN());
   DFF_X1 \o_values_reg[55][8]  (.D(o_values[8]), .CK(n_0_112), .Q(
      \o_values[55] [8]), .QN());
   DFF_X1 \o_values_reg[55][7]  (.D(o_values[7]), .CK(n_0_112), .Q(
      \o_values[55] [7]), .QN());
   DFF_X1 \o_values_reg[55][6]  (.D(o_values[6]), .CK(n_0_112), .Q(
      \o_values[55] [6]), .QN());
   DFF_X1 \o_values_reg[55][5]  (.D(o_values[5]), .CK(n_0_112), .Q(
      \o_values[55] [5]), .QN());
   DFF_X1 \o_values_reg[55][4]  (.D(o_values[4]), .CK(n_0_112), .Q(
      \o_values[55] [4]), .QN());
   DFF_X1 \o_values_reg[55][3]  (.D(o_values[3]), .CK(n_0_112), .Q(
      \o_values[55] [3]), .QN());
   DFF_X1 \o_values_reg[55][2]  (.D(o_values[2]), .CK(n_0_112), .Q(
      \o_values[55] [2]), .QN());
   DFF_X1 \o_values_reg[55][1]  (.D(o_values[1]), .CK(n_0_112), .Q(
      \o_values[55] [1]), .QN());
   DFF_X1 \o_values_reg[55][0]  (.D(o_values[0]), .CK(n_0_112), .Q(
      \o_values[55] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[54]_reg  (.CK(clk), .E(n_0_29), .SE(1'b0), 
      .GCK(n_0_113));
   DFF_X1 \o_values_reg[54][15]  (.D(o_values[15]), .CK(n_0_113), .Q(
      \o_values[54] [15]), .QN());
   DFF_X1 \o_values_reg[54][14]  (.D(o_values[14]), .CK(n_0_113), .Q(
      \o_values[54] [14]), .QN());
   DFF_X1 \o_values_reg[54][13]  (.D(o_values[13]), .CK(n_0_113), .Q(
      \o_values[54] [13]), .QN());
   DFF_X1 \o_values_reg[54][12]  (.D(o_values[12]), .CK(n_0_113), .Q(
      \o_values[54] [12]), .QN());
   DFF_X1 \o_values_reg[54][11]  (.D(o_values[11]), .CK(n_0_113), .Q(
      \o_values[54] [11]), .QN());
   DFF_X1 \o_values_reg[54][10]  (.D(o_values[10]), .CK(n_0_113), .Q(
      \o_values[54] [10]), .QN());
   DFF_X1 \o_values_reg[54][9]  (.D(o_values[9]), .CK(n_0_113), .Q(
      \o_values[54] [9]), .QN());
   DFF_X1 \o_values_reg[54][8]  (.D(o_values[8]), .CK(n_0_113), .Q(
      \o_values[54] [8]), .QN());
   DFF_X1 \o_values_reg[54][7]  (.D(o_values[7]), .CK(n_0_113), .Q(
      \o_values[54] [7]), .QN());
   DFF_X1 \o_values_reg[54][6]  (.D(o_values[6]), .CK(n_0_113), .Q(
      \o_values[54] [6]), .QN());
   DFF_X1 \o_values_reg[54][5]  (.D(o_values[5]), .CK(n_0_113), .Q(
      \o_values[54] [5]), .QN());
   DFF_X1 \o_values_reg[54][4]  (.D(o_values[4]), .CK(n_0_113), .Q(
      \o_values[54] [4]), .QN());
   DFF_X1 \o_values_reg[54][3]  (.D(o_values[3]), .CK(n_0_113), .Q(
      \o_values[54] [3]), .QN());
   DFF_X1 \o_values_reg[54][2]  (.D(o_values[2]), .CK(n_0_113), .Q(
      \o_values[54] [2]), .QN());
   DFF_X1 \o_values_reg[54][1]  (.D(o_values[1]), .CK(n_0_113), .Q(
      \o_values[54] [1]), .QN());
   DFF_X1 \o_values_reg[54][0]  (.D(o_values[0]), .CK(n_0_113), .Q(
      \o_values[54] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[53]_reg  (.CK(clk), .E(n_0_30), .SE(1'b0), 
      .GCK(n_0_114));
   DFF_X1 \o_values_reg[53][15]  (.D(o_values[15]), .CK(n_0_114), .Q(
      \o_values[53] [15]), .QN());
   DFF_X1 \o_values_reg[53][14]  (.D(o_values[14]), .CK(n_0_114), .Q(
      \o_values[53] [14]), .QN());
   DFF_X1 \o_values_reg[53][13]  (.D(o_values[13]), .CK(n_0_114), .Q(
      \o_values[53] [13]), .QN());
   DFF_X1 \o_values_reg[53][12]  (.D(o_values[12]), .CK(n_0_114), .Q(
      \o_values[53] [12]), .QN());
   DFF_X1 \o_values_reg[53][11]  (.D(o_values[11]), .CK(n_0_114), .Q(
      \o_values[53] [11]), .QN());
   DFF_X1 \o_values_reg[53][10]  (.D(o_values[10]), .CK(n_0_114), .Q(
      \o_values[53] [10]), .QN());
   DFF_X1 \o_values_reg[53][9]  (.D(o_values[9]), .CK(n_0_114), .Q(
      \o_values[53] [9]), .QN());
   DFF_X1 \o_values_reg[53][8]  (.D(o_values[8]), .CK(n_0_114), .Q(
      \o_values[53] [8]), .QN());
   DFF_X1 \o_values_reg[53][7]  (.D(o_values[7]), .CK(n_0_114), .Q(
      \o_values[53] [7]), .QN());
   DFF_X1 \o_values_reg[53][6]  (.D(o_values[6]), .CK(n_0_114), .Q(
      \o_values[53] [6]), .QN());
   DFF_X1 \o_values_reg[53][5]  (.D(o_values[5]), .CK(n_0_114), .Q(
      \o_values[53] [5]), .QN());
   DFF_X1 \o_values_reg[53][4]  (.D(o_values[4]), .CK(n_0_114), .Q(
      \o_values[53] [4]), .QN());
   DFF_X1 \o_values_reg[53][3]  (.D(o_values[3]), .CK(n_0_114), .Q(
      \o_values[53] [3]), .QN());
   DFF_X1 \o_values_reg[53][2]  (.D(o_values[2]), .CK(n_0_114), .Q(
      \o_values[53] [2]), .QN());
   DFF_X1 \o_values_reg[53][1]  (.D(o_values[1]), .CK(n_0_114), .Q(
      \o_values[53] [1]), .QN());
   DFF_X1 \o_values_reg[53][0]  (.D(o_values[0]), .CK(n_0_114), .Q(
      \o_values[53] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[52]_reg  (.CK(clk), .E(n_0_31), .SE(1'b0), 
      .GCK(n_0_115));
   DFF_X1 \o_values_reg[52][15]  (.D(o_values[15]), .CK(n_0_115), .Q(
      \o_values[52] [15]), .QN());
   DFF_X1 \o_values_reg[52][14]  (.D(o_values[14]), .CK(n_0_115), .Q(
      \o_values[52] [14]), .QN());
   DFF_X1 \o_values_reg[52][13]  (.D(o_values[13]), .CK(n_0_115), .Q(
      \o_values[52] [13]), .QN());
   DFF_X1 \o_values_reg[52][12]  (.D(o_values[12]), .CK(n_0_115), .Q(
      \o_values[52] [12]), .QN());
   DFF_X1 \o_values_reg[52][11]  (.D(o_values[11]), .CK(n_0_115), .Q(
      \o_values[52] [11]), .QN());
   DFF_X1 \o_values_reg[52][10]  (.D(o_values[10]), .CK(n_0_115), .Q(
      \o_values[52] [10]), .QN());
   DFF_X1 \o_values_reg[52][9]  (.D(o_values[9]), .CK(n_0_115), .Q(
      \o_values[52] [9]), .QN());
   DFF_X1 \o_values_reg[52][8]  (.D(o_values[8]), .CK(n_0_115), .Q(
      \o_values[52] [8]), .QN());
   DFF_X1 \o_values_reg[52][7]  (.D(o_values[7]), .CK(n_0_115), .Q(
      \o_values[52] [7]), .QN());
   DFF_X1 \o_values_reg[52][6]  (.D(o_values[6]), .CK(n_0_115), .Q(
      \o_values[52] [6]), .QN());
   DFF_X1 \o_values_reg[52][5]  (.D(o_values[5]), .CK(n_0_115), .Q(
      \o_values[52] [5]), .QN());
   DFF_X1 \o_values_reg[52][4]  (.D(o_values[4]), .CK(n_0_115), .Q(
      \o_values[52] [4]), .QN());
   DFF_X1 \o_values_reg[52][3]  (.D(o_values[3]), .CK(n_0_115), .Q(
      \o_values[52] [3]), .QN());
   DFF_X1 \o_values_reg[52][2]  (.D(o_values[2]), .CK(n_0_115), .Q(
      \o_values[52] [2]), .QN());
   DFF_X1 \o_values_reg[52][1]  (.D(o_values[1]), .CK(n_0_115), .Q(
      \o_values[52] [1]), .QN());
   DFF_X1 \o_values_reg[52][0]  (.D(o_values[0]), .CK(n_0_115), .Q(
      \o_values[52] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[51]_reg  (.CK(clk), .E(n_0_32), .SE(1'b0), 
      .GCK(n_0_116));
   DFF_X1 \o_values_reg[51][15]  (.D(o_values[15]), .CK(n_0_116), .Q(
      \o_values[51] [15]), .QN());
   DFF_X1 \o_values_reg[51][14]  (.D(o_values[14]), .CK(n_0_116), .Q(
      \o_values[51] [14]), .QN());
   DFF_X1 \o_values_reg[51][13]  (.D(o_values[13]), .CK(n_0_116), .Q(
      \o_values[51] [13]), .QN());
   DFF_X1 \o_values_reg[51][12]  (.D(o_values[12]), .CK(n_0_116), .Q(
      \o_values[51] [12]), .QN());
   DFF_X1 \o_values_reg[51][11]  (.D(o_values[11]), .CK(n_0_116), .Q(
      \o_values[51] [11]), .QN());
   DFF_X1 \o_values_reg[51][10]  (.D(o_values[10]), .CK(n_0_116), .Q(
      \o_values[51] [10]), .QN());
   DFF_X1 \o_values_reg[51][9]  (.D(o_values[9]), .CK(n_0_116), .Q(
      \o_values[51] [9]), .QN());
   DFF_X1 \o_values_reg[51][8]  (.D(o_values[8]), .CK(n_0_116), .Q(
      \o_values[51] [8]), .QN());
   DFF_X1 \o_values_reg[51][7]  (.D(o_values[7]), .CK(n_0_116), .Q(
      \o_values[51] [7]), .QN());
   DFF_X1 \o_values_reg[51][6]  (.D(o_values[6]), .CK(n_0_116), .Q(
      \o_values[51] [6]), .QN());
   DFF_X1 \o_values_reg[51][5]  (.D(o_values[5]), .CK(n_0_116), .Q(
      \o_values[51] [5]), .QN());
   DFF_X1 \o_values_reg[51][4]  (.D(o_values[4]), .CK(n_0_116), .Q(
      \o_values[51] [4]), .QN());
   DFF_X1 \o_values_reg[51][3]  (.D(o_values[3]), .CK(n_0_116), .Q(
      \o_values[51] [3]), .QN());
   DFF_X1 \o_values_reg[51][2]  (.D(o_values[2]), .CK(n_0_116), .Q(
      \o_values[51] [2]), .QN());
   DFF_X1 \o_values_reg[51][1]  (.D(o_values[1]), .CK(n_0_116), .Q(
      \o_values[51] [1]), .QN());
   DFF_X1 \o_values_reg[51][0]  (.D(o_values[0]), .CK(n_0_116), .Q(
      \o_values[51] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[50]_reg  (.CK(clk), .E(n_0_33), .SE(1'b0), 
      .GCK(n_0_117));
   DFF_X1 \o_values_reg[50][15]  (.D(o_values[15]), .CK(n_0_117), .Q(
      \o_values[50] [15]), .QN());
   DFF_X1 \o_values_reg[50][14]  (.D(o_values[14]), .CK(n_0_117), .Q(
      \o_values[50] [14]), .QN());
   DFF_X1 \o_values_reg[50][13]  (.D(o_values[13]), .CK(n_0_117), .Q(
      \o_values[50] [13]), .QN());
   DFF_X1 \o_values_reg[50][12]  (.D(o_values[12]), .CK(n_0_117), .Q(
      \o_values[50] [12]), .QN());
   DFF_X1 \o_values_reg[50][11]  (.D(o_values[11]), .CK(n_0_117), .Q(
      \o_values[50] [11]), .QN());
   DFF_X1 \o_values_reg[50][10]  (.D(o_values[10]), .CK(n_0_117), .Q(
      \o_values[50] [10]), .QN());
   DFF_X1 \o_values_reg[50][9]  (.D(o_values[9]), .CK(n_0_117), .Q(
      \o_values[50] [9]), .QN());
   DFF_X1 \o_values_reg[50][8]  (.D(o_values[8]), .CK(n_0_117), .Q(
      \o_values[50] [8]), .QN());
   DFF_X1 \o_values_reg[50][7]  (.D(o_values[7]), .CK(n_0_117), .Q(
      \o_values[50] [7]), .QN());
   DFF_X1 \o_values_reg[50][6]  (.D(o_values[6]), .CK(n_0_117), .Q(
      \o_values[50] [6]), .QN());
   DFF_X1 \o_values_reg[50][5]  (.D(o_values[5]), .CK(n_0_117), .Q(
      \o_values[50] [5]), .QN());
   DFF_X1 \o_values_reg[50][4]  (.D(o_values[4]), .CK(n_0_117), .Q(
      \o_values[50] [4]), .QN());
   DFF_X1 \o_values_reg[50][3]  (.D(o_values[3]), .CK(n_0_117), .Q(
      \o_values[50] [3]), .QN());
   DFF_X1 \o_values_reg[50][2]  (.D(o_values[2]), .CK(n_0_117), .Q(
      \o_values[50] [2]), .QN());
   DFF_X1 \o_values_reg[50][1]  (.D(o_values[1]), .CK(n_0_117), .Q(
      \o_values[50] [1]), .QN());
   DFF_X1 \o_values_reg[50][0]  (.D(o_values[0]), .CK(n_0_117), .Q(
      \o_values[50] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[49]_reg  (.CK(clk), .E(n_0_34), .SE(1'b0), 
      .GCK(n_0_118));
   DFF_X1 \o_values_reg[49][15]  (.D(o_values[15]), .CK(n_0_118), .Q(
      \o_values[49] [15]), .QN());
   DFF_X1 \o_values_reg[49][14]  (.D(o_values[14]), .CK(n_0_118), .Q(
      \o_values[49] [14]), .QN());
   DFF_X1 \o_values_reg[49][13]  (.D(o_values[13]), .CK(n_0_118), .Q(
      \o_values[49] [13]), .QN());
   DFF_X1 \o_values_reg[49][12]  (.D(o_values[12]), .CK(n_0_118), .Q(
      \o_values[49] [12]), .QN());
   DFF_X1 \o_values_reg[49][11]  (.D(o_values[11]), .CK(n_0_118), .Q(
      \o_values[49] [11]), .QN());
   DFF_X1 \o_values_reg[49][10]  (.D(o_values[10]), .CK(n_0_118), .Q(
      \o_values[49] [10]), .QN());
   DFF_X1 \o_values_reg[49][9]  (.D(o_values[9]), .CK(n_0_118), .Q(
      \o_values[49] [9]), .QN());
   DFF_X1 \o_values_reg[49][8]  (.D(o_values[8]), .CK(n_0_118), .Q(
      \o_values[49] [8]), .QN());
   DFF_X1 \o_values_reg[49][7]  (.D(o_values[7]), .CK(n_0_118), .Q(
      \o_values[49] [7]), .QN());
   DFF_X1 \o_values_reg[49][6]  (.D(o_values[6]), .CK(n_0_118), .Q(
      \o_values[49] [6]), .QN());
   DFF_X1 \o_values_reg[49][5]  (.D(o_values[5]), .CK(n_0_118), .Q(
      \o_values[49] [5]), .QN());
   DFF_X1 \o_values_reg[49][4]  (.D(o_values[4]), .CK(n_0_118), .Q(
      \o_values[49] [4]), .QN());
   DFF_X1 \o_values_reg[49][3]  (.D(o_values[3]), .CK(n_0_118), .Q(
      \o_values[49] [3]), .QN());
   DFF_X1 \o_values_reg[49][2]  (.D(o_values[2]), .CK(n_0_118), .Q(
      \o_values[49] [2]), .QN());
   DFF_X1 \o_values_reg[49][1]  (.D(o_values[1]), .CK(n_0_118), .Q(
      \o_values[49] [1]), .QN());
   DFF_X1 \o_values_reg[49][0]  (.D(o_values[0]), .CK(n_0_118), .Q(
      \o_values[49] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[48]_reg  (.CK(clk), .E(n_0_35), .SE(1'b0), 
      .GCK(n_0_119));
   DFF_X1 \o_values_reg[48][15]  (.D(o_values[15]), .CK(n_0_119), .Q(
      \o_values[48] [15]), .QN());
   DFF_X1 \o_values_reg[48][14]  (.D(o_values[14]), .CK(n_0_119), .Q(
      \o_values[48] [14]), .QN());
   DFF_X1 \o_values_reg[48][13]  (.D(o_values[13]), .CK(n_0_119), .Q(
      \o_values[48] [13]), .QN());
   DFF_X1 \o_values_reg[48][12]  (.D(o_values[12]), .CK(n_0_119), .Q(
      \o_values[48] [12]), .QN());
   DFF_X1 \o_values_reg[48][11]  (.D(o_values[11]), .CK(n_0_119), .Q(
      \o_values[48] [11]), .QN());
   DFF_X1 \o_values_reg[48][10]  (.D(o_values[10]), .CK(n_0_119), .Q(
      \o_values[48] [10]), .QN());
   DFF_X1 \o_values_reg[48][9]  (.D(o_values[9]), .CK(n_0_119), .Q(
      \o_values[48] [9]), .QN());
   DFF_X1 \o_values_reg[48][8]  (.D(o_values[8]), .CK(n_0_119), .Q(
      \o_values[48] [8]), .QN());
   DFF_X1 \o_values_reg[48][7]  (.D(o_values[7]), .CK(n_0_119), .Q(
      \o_values[48] [7]), .QN());
   DFF_X1 \o_values_reg[48][6]  (.D(o_values[6]), .CK(n_0_119), .Q(
      \o_values[48] [6]), .QN());
   DFF_X1 \o_values_reg[48][5]  (.D(o_values[5]), .CK(n_0_119), .Q(
      \o_values[48] [5]), .QN());
   DFF_X1 \o_values_reg[48][4]  (.D(o_values[4]), .CK(n_0_119), .Q(
      \o_values[48] [4]), .QN());
   DFF_X1 \o_values_reg[48][3]  (.D(o_values[3]), .CK(n_0_119), .Q(
      \o_values[48] [3]), .QN());
   DFF_X1 \o_values_reg[48][2]  (.D(o_values[2]), .CK(n_0_119), .Q(
      \o_values[48] [2]), .QN());
   DFF_X1 \o_values_reg[48][1]  (.D(o_values[1]), .CK(n_0_119), .Q(
      \o_values[48] [1]), .QN());
   DFF_X1 \o_values_reg[48][0]  (.D(o_values[0]), .CK(n_0_119), .Q(
      \o_values[48] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[47]_reg  (.CK(clk), .E(n_0_36), .SE(1'b0), 
      .GCK(n_0_120));
   DFF_X1 \o_values_reg[47][15]  (.D(o_values[15]), .CK(n_0_120), .Q(
      \o_values[47] [15]), .QN());
   DFF_X1 \o_values_reg[47][14]  (.D(o_values[14]), .CK(n_0_120), .Q(
      \o_values[47] [14]), .QN());
   DFF_X1 \o_values_reg[47][13]  (.D(o_values[13]), .CK(n_0_120), .Q(
      \o_values[47] [13]), .QN());
   DFF_X1 \o_values_reg[47][12]  (.D(o_values[12]), .CK(n_0_120), .Q(
      \o_values[47] [12]), .QN());
   DFF_X1 \o_values_reg[47][11]  (.D(o_values[11]), .CK(n_0_120), .Q(
      \o_values[47] [11]), .QN());
   DFF_X1 \o_values_reg[47][10]  (.D(o_values[10]), .CK(n_0_120), .Q(
      \o_values[47] [10]), .QN());
   DFF_X1 \o_values_reg[47][9]  (.D(o_values[9]), .CK(n_0_120), .Q(
      \o_values[47] [9]), .QN());
   DFF_X1 \o_values_reg[47][8]  (.D(o_values[8]), .CK(n_0_120), .Q(
      \o_values[47] [8]), .QN());
   DFF_X1 \o_values_reg[47][7]  (.D(o_values[7]), .CK(n_0_120), .Q(
      \o_values[47] [7]), .QN());
   DFF_X1 \o_values_reg[47][6]  (.D(o_values[6]), .CK(n_0_120), .Q(
      \o_values[47] [6]), .QN());
   DFF_X1 \o_values_reg[47][5]  (.D(o_values[5]), .CK(n_0_120), .Q(
      \o_values[47] [5]), .QN());
   DFF_X1 \o_values_reg[47][4]  (.D(o_values[4]), .CK(n_0_120), .Q(
      \o_values[47] [4]), .QN());
   DFF_X1 \o_values_reg[47][3]  (.D(o_values[3]), .CK(n_0_120), .Q(
      \o_values[47] [3]), .QN());
   DFF_X1 \o_values_reg[47][2]  (.D(o_values[2]), .CK(n_0_120), .Q(
      \o_values[47] [2]), .QN());
   DFF_X1 \o_values_reg[47][1]  (.D(o_values[1]), .CK(n_0_120), .Q(
      \o_values[47] [1]), .QN());
   DFF_X1 \o_values_reg[47][0]  (.D(o_values[0]), .CK(n_0_120), .Q(
      \o_values[47] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[46]_reg  (.CK(clk), .E(n_0_37), .SE(1'b0), 
      .GCK(n_0_121));
   DFF_X1 \o_values_reg[46][15]  (.D(o_values[15]), .CK(n_0_121), .Q(
      \o_values[46] [15]), .QN());
   DFF_X1 \o_values_reg[46][14]  (.D(o_values[14]), .CK(n_0_121), .Q(
      \o_values[46] [14]), .QN());
   DFF_X1 \o_values_reg[46][13]  (.D(o_values[13]), .CK(n_0_121), .Q(
      \o_values[46] [13]), .QN());
   DFF_X1 \o_values_reg[46][12]  (.D(o_values[12]), .CK(n_0_121), .Q(
      \o_values[46] [12]), .QN());
   DFF_X1 \o_values_reg[46][11]  (.D(o_values[11]), .CK(n_0_121), .Q(
      \o_values[46] [11]), .QN());
   DFF_X1 \o_values_reg[46][10]  (.D(o_values[10]), .CK(n_0_121), .Q(
      \o_values[46] [10]), .QN());
   DFF_X1 \o_values_reg[46][9]  (.D(o_values[9]), .CK(n_0_121), .Q(
      \o_values[46] [9]), .QN());
   DFF_X1 \o_values_reg[46][8]  (.D(o_values[8]), .CK(n_0_121), .Q(
      \o_values[46] [8]), .QN());
   DFF_X1 \o_values_reg[46][7]  (.D(o_values[7]), .CK(n_0_121), .Q(
      \o_values[46] [7]), .QN());
   DFF_X1 \o_values_reg[46][6]  (.D(o_values[6]), .CK(n_0_121), .Q(
      \o_values[46] [6]), .QN());
   DFF_X1 \o_values_reg[46][5]  (.D(o_values[5]), .CK(n_0_121), .Q(
      \o_values[46] [5]), .QN());
   DFF_X1 \o_values_reg[46][4]  (.D(o_values[4]), .CK(n_0_121), .Q(
      \o_values[46] [4]), .QN());
   DFF_X1 \o_values_reg[46][3]  (.D(o_values[3]), .CK(n_0_121), .Q(
      \o_values[46] [3]), .QN());
   DFF_X1 \o_values_reg[46][2]  (.D(o_values[2]), .CK(n_0_121), .Q(
      \o_values[46] [2]), .QN());
   DFF_X1 \o_values_reg[46][1]  (.D(o_values[1]), .CK(n_0_121), .Q(
      \o_values[46] [1]), .QN());
   DFF_X1 \o_values_reg[46][0]  (.D(o_values[0]), .CK(n_0_121), .Q(
      \o_values[46] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[45]_reg  (.CK(clk), .E(n_0_38), .SE(1'b0), 
      .GCK(n_0_122));
   DFF_X1 \o_values_reg[45][15]  (.D(o_values[15]), .CK(n_0_122), .Q(
      \o_values[45] [15]), .QN());
   DFF_X1 \o_values_reg[45][14]  (.D(o_values[14]), .CK(n_0_122), .Q(
      \o_values[45] [14]), .QN());
   DFF_X1 \o_values_reg[45][13]  (.D(o_values[13]), .CK(n_0_122), .Q(
      \o_values[45] [13]), .QN());
   DFF_X1 \o_values_reg[45][12]  (.D(o_values[12]), .CK(n_0_122), .Q(
      \o_values[45] [12]), .QN());
   DFF_X1 \o_values_reg[45][11]  (.D(o_values[11]), .CK(n_0_122), .Q(
      \o_values[45] [11]), .QN());
   DFF_X1 \o_values_reg[45][10]  (.D(o_values[10]), .CK(n_0_122), .Q(
      \o_values[45] [10]), .QN());
   DFF_X1 \o_values_reg[45][9]  (.D(o_values[9]), .CK(n_0_122), .Q(
      \o_values[45] [9]), .QN());
   DFF_X1 \o_values_reg[45][8]  (.D(o_values[8]), .CK(n_0_122), .Q(
      \o_values[45] [8]), .QN());
   DFF_X1 \o_values_reg[45][7]  (.D(o_values[7]), .CK(n_0_122), .Q(
      \o_values[45] [7]), .QN());
   DFF_X1 \o_values_reg[45][6]  (.D(o_values[6]), .CK(n_0_122), .Q(
      \o_values[45] [6]), .QN());
   DFF_X1 \o_values_reg[45][5]  (.D(o_values[5]), .CK(n_0_122), .Q(
      \o_values[45] [5]), .QN());
   DFF_X1 \o_values_reg[45][4]  (.D(o_values[4]), .CK(n_0_122), .Q(
      \o_values[45] [4]), .QN());
   DFF_X1 \o_values_reg[45][3]  (.D(o_values[3]), .CK(n_0_122), .Q(
      \o_values[45] [3]), .QN());
   DFF_X1 \o_values_reg[45][2]  (.D(o_values[2]), .CK(n_0_122), .Q(
      \o_values[45] [2]), .QN());
   DFF_X1 \o_values_reg[45][1]  (.D(o_values[1]), .CK(n_0_122), .Q(
      \o_values[45] [1]), .QN());
   DFF_X1 \o_values_reg[45][0]  (.D(o_values[0]), .CK(n_0_122), .Q(
      \o_values[45] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[44]_reg  (.CK(clk), .E(n_0_39), .SE(1'b0), 
      .GCK(n_0_123));
   DFF_X1 \o_values_reg[44][15]  (.D(o_values[15]), .CK(n_0_123), .Q(
      \o_values[44] [15]), .QN());
   DFF_X1 \o_values_reg[44][14]  (.D(o_values[14]), .CK(n_0_123), .Q(
      \o_values[44] [14]), .QN());
   DFF_X1 \o_values_reg[44][13]  (.D(o_values[13]), .CK(n_0_123), .Q(
      \o_values[44] [13]), .QN());
   DFF_X1 \o_values_reg[44][12]  (.D(o_values[12]), .CK(n_0_123), .Q(
      \o_values[44] [12]), .QN());
   DFF_X1 \o_values_reg[44][11]  (.D(o_values[11]), .CK(n_0_123), .Q(
      \o_values[44] [11]), .QN());
   DFF_X1 \o_values_reg[44][10]  (.D(o_values[10]), .CK(n_0_123), .Q(
      \o_values[44] [10]), .QN());
   DFF_X1 \o_values_reg[44][9]  (.D(o_values[9]), .CK(n_0_123), .Q(
      \o_values[44] [9]), .QN());
   DFF_X1 \o_values_reg[44][8]  (.D(o_values[8]), .CK(n_0_123), .Q(
      \o_values[44] [8]), .QN());
   DFF_X1 \o_values_reg[44][7]  (.D(o_values[7]), .CK(n_0_123), .Q(
      \o_values[44] [7]), .QN());
   DFF_X1 \o_values_reg[44][6]  (.D(o_values[6]), .CK(n_0_123), .Q(
      \o_values[44] [6]), .QN());
   DFF_X1 \o_values_reg[44][5]  (.D(o_values[5]), .CK(n_0_123), .Q(
      \o_values[44] [5]), .QN());
   DFF_X1 \o_values_reg[44][4]  (.D(o_values[4]), .CK(n_0_123), .Q(
      \o_values[44] [4]), .QN());
   DFF_X1 \o_values_reg[44][3]  (.D(o_values[3]), .CK(n_0_123), .Q(
      \o_values[44] [3]), .QN());
   DFF_X1 \o_values_reg[44][2]  (.D(o_values[2]), .CK(n_0_123), .Q(
      \o_values[44] [2]), .QN());
   DFF_X1 \o_values_reg[44][1]  (.D(o_values[1]), .CK(n_0_123), .Q(
      \o_values[44] [1]), .QN());
   DFF_X1 \o_values_reg[44][0]  (.D(o_values[0]), .CK(n_0_123), .Q(
      \o_values[44] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[43]_reg  (.CK(clk), .E(n_0_40), .SE(1'b0), 
      .GCK(n_0_124));
   DFF_X1 \o_values_reg[43][15]  (.D(o_values[15]), .CK(n_0_124), .Q(
      \o_values[43] [15]), .QN());
   DFF_X1 \o_values_reg[43][14]  (.D(o_values[14]), .CK(n_0_124), .Q(
      \o_values[43] [14]), .QN());
   DFF_X1 \o_values_reg[43][13]  (.D(o_values[13]), .CK(n_0_124), .Q(
      \o_values[43] [13]), .QN());
   DFF_X1 \o_values_reg[43][12]  (.D(o_values[12]), .CK(n_0_124), .Q(
      \o_values[43] [12]), .QN());
   DFF_X1 \o_values_reg[43][11]  (.D(o_values[11]), .CK(n_0_124), .Q(
      \o_values[43] [11]), .QN());
   DFF_X1 \o_values_reg[43][10]  (.D(o_values[10]), .CK(n_0_124), .Q(
      \o_values[43] [10]), .QN());
   DFF_X1 \o_values_reg[43][9]  (.D(o_values[9]), .CK(n_0_124), .Q(
      \o_values[43] [9]), .QN());
   DFF_X1 \o_values_reg[43][8]  (.D(o_values[8]), .CK(n_0_124), .Q(
      \o_values[43] [8]), .QN());
   DFF_X1 \o_values_reg[43][7]  (.D(o_values[7]), .CK(n_0_124), .Q(
      \o_values[43] [7]), .QN());
   DFF_X1 \o_values_reg[43][6]  (.D(o_values[6]), .CK(n_0_124), .Q(
      \o_values[43] [6]), .QN());
   DFF_X1 \o_values_reg[43][5]  (.D(o_values[5]), .CK(n_0_124), .Q(
      \o_values[43] [5]), .QN());
   DFF_X1 \o_values_reg[43][4]  (.D(o_values[4]), .CK(n_0_124), .Q(
      \o_values[43] [4]), .QN());
   DFF_X1 \o_values_reg[43][3]  (.D(o_values[3]), .CK(n_0_124), .Q(
      \o_values[43] [3]), .QN());
   DFF_X1 \o_values_reg[43][2]  (.D(o_values[2]), .CK(n_0_124), .Q(
      \o_values[43] [2]), .QN());
   DFF_X1 \o_values_reg[43][1]  (.D(o_values[1]), .CK(n_0_124), .Q(
      \o_values[43] [1]), .QN());
   DFF_X1 \o_values_reg[43][0]  (.D(o_values[0]), .CK(n_0_124), .Q(
      \o_values[43] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[42]_reg  (.CK(clk), .E(n_0_41), .SE(1'b0), 
      .GCK(n_0_125));
   DFF_X1 \o_values_reg[42][15]  (.D(o_values[15]), .CK(n_0_125), .Q(
      \o_values[42] [15]), .QN());
   DFF_X1 \o_values_reg[42][14]  (.D(o_values[14]), .CK(n_0_125), .Q(
      \o_values[42] [14]), .QN());
   DFF_X1 \o_values_reg[42][13]  (.D(o_values[13]), .CK(n_0_125), .Q(
      \o_values[42] [13]), .QN());
   DFF_X1 \o_values_reg[42][12]  (.D(o_values[12]), .CK(n_0_125), .Q(
      \o_values[42] [12]), .QN());
   DFF_X1 \o_values_reg[42][11]  (.D(o_values[11]), .CK(n_0_125), .Q(
      \o_values[42] [11]), .QN());
   DFF_X1 \o_values_reg[42][10]  (.D(o_values[10]), .CK(n_0_125), .Q(
      \o_values[42] [10]), .QN());
   DFF_X1 \o_values_reg[42][9]  (.D(o_values[9]), .CK(n_0_125), .Q(
      \o_values[42] [9]), .QN());
   DFF_X1 \o_values_reg[42][8]  (.D(o_values[8]), .CK(n_0_125), .Q(
      \o_values[42] [8]), .QN());
   DFF_X1 \o_values_reg[42][7]  (.D(o_values[7]), .CK(n_0_125), .Q(
      \o_values[42] [7]), .QN());
   DFF_X1 \o_values_reg[42][6]  (.D(o_values[6]), .CK(n_0_125), .Q(
      \o_values[42] [6]), .QN());
   DFF_X1 \o_values_reg[42][5]  (.D(o_values[5]), .CK(n_0_125), .Q(
      \o_values[42] [5]), .QN());
   DFF_X1 \o_values_reg[42][4]  (.D(o_values[4]), .CK(n_0_125), .Q(
      \o_values[42] [4]), .QN());
   DFF_X1 \o_values_reg[42][3]  (.D(o_values[3]), .CK(n_0_125), .Q(
      \o_values[42] [3]), .QN());
   DFF_X1 \o_values_reg[42][2]  (.D(o_values[2]), .CK(n_0_125), .Q(
      \o_values[42] [2]), .QN());
   DFF_X1 \o_values_reg[42][1]  (.D(o_values[1]), .CK(n_0_125), .Q(
      \o_values[42] [1]), .QN());
   DFF_X1 \o_values_reg[42][0]  (.D(o_values[0]), .CK(n_0_125), .Q(
      \o_values[42] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[41]_reg  (.CK(clk), .E(n_0_42), .SE(1'b0), 
      .GCK(n_0_126));
   DFF_X1 \o_values_reg[41][15]  (.D(o_values[15]), .CK(n_0_126), .Q(
      \o_values[41] [15]), .QN());
   DFF_X1 \o_values_reg[41][14]  (.D(o_values[14]), .CK(n_0_126), .Q(
      \o_values[41] [14]), .QN());
   DFF_X1 \o_values_reg[41][13]  (.D(o_values[13]), .CK(n_0_126), .Q(
      \o_values[41] [13]), .QN());
   DFF_X1 \o_values_reg[41][12]  (.D(o_values[12]), .CK(n_0_126), .Q(
      \o_values[41] [12]), .QN());
   DFF_X1 \o_values_reg[41][11]  (.D(o_values[11]), .CK(n_0_126), .Q(
      \o_values[41] [11]), .QN());
   DFF_X1 \o_values_reg[41][10]  (.D(o_values[10]), .CK(n_0_126), .Q(
      \o_values[41] [10]), .QN());
   DFF_X1 \o_values_reg[41][9]  (.D(o_values[9]), .CK(n_0_126), .Q(
      \o_values[41] [9]), .QN());
   DFF_X1 \o_values_reg[41][8]  (.D(o_values[8]), .CK(n_0_126), .Q(
      \o_values[41] [8]), .QN());
   DFF_X1 \o_values_reg[41][7]  (.D(o_values[7]), .CK(n_0_126), .Q(
      \o_values[41] [7]), .QN());
   DFF_X1 \o_values_reg[41][6]  (.D(o_values[6]), .CK(n_0_126), .Q(
      \o_values[41] [6]), .QN());
   DFF_X1 \o_values_reg[41][5]  (.D(o_values[5]), .CK(n_0_126), .Q(
      \o_values[41] [5]), .QN());
   DFF_X1 \o_values_reg[41][4]  (.D(o_values[4]), .CK(n_0_126), .Q(
      \o_values[41] [4]), .QN());
   DFF_X1 \o_values_reg[41][3]  (.D(o_values[3]), .CK(n_0_126), .Q(
      \o_values[41] [3]), .QN());
   DFF_X1 \o_values_reg[41][2]  (.D(o_values[2]), .CK(n_0_126), .Q(
      \o_values[41] [2]), .QN());
   DFF_X1 \o_values_reg[41][1]  (.D(o_values[1]), .CK(n_0_126), .Q(
      \o_values[41] [1]), .QN());
   DFF_X1 \o_values_reg[41][0]  (.D(o_values[0]), .CK(n_0_126), .Q(
      \o_values[41] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[40]_reg  (.CK(clk), .E(n_0_43), .SE(1'b0), 
      .GCK(n_0_127));
   DFF_X1 \o_values_reg[40][15]  (.D(o_values[15]), .CK(n_0_127), .Q(
      \o_values[40] [15]), .QN());
   DFF_X1 \o_values_reg[40][14]  (.D(o_values[14]), .CK(n_0_127), .Q(
      \o_values[40] [14]), .QN());
   DFF_X1 \o_values_reg[40][13]  (.D(o_values[13]), .CK(n_0_127), .Q(
      \o_values[40] [13]), .QN());
   DFF_X1 \o_values_reg[40][12]  (.D(o_values[12]), .CK(n_0_127), .Q(
      \o_values[40] [12]), .QN());
   DFF_X1 \o_values_reg[40][11]  (.D(o_values[11]), .CK(n_0_127), .Q(
      \o_values[40] [11]), .QN());
   DFF_X1 \o_values_reg[40][10]  (.D(o_values[10]), .CK(n_0_127), .Q(
      \o_values[40] [10]), .QN());
   DFF_X1 \o_values_reg[40][9]  (.D(o_values[9]), .CK(n_0_127), .Q(
      \o_values[40] [9]), .QN());
   DFF_X1 \o_values_reg[40][8]  (.D(o_values[8]), .CK(n_0_127), .Q(
      \o_values[40] [8]), .QN());
   DFF_X1 \o_values_reg[40][7]  (.D(o_values[7]), .CK(n_0_127), .Q(
      \o_values[40] [7]), .QN());
   DFF_X1 \o_values_reg[40][6]  (.D(o_values[6]), .CK(n_0_127), .Q(
      \o_values[40] [6]), .QN());
   DFF_X1 \o_values_reg[40][5]  (.D(o_values[5]), .CK(n_0_127), .Q(
      \o_values[40] [5]), .QN());
   DFF_X1 \o_values_reg[40][4]  (.D(o_values[4]), .CK(n_0_127), .Q(
      \o_values[40] [4]), .QN());
   DFF_X1 \o_values_reg[40][3]  (.D(o_values[3]), .CK(n_0_127), .Q(
      \o_values[40] [3]), .QN());
   DFF_X1 \o_values_reg[40][2]  (.D(o_values[2]), .CK(n_0_127), .Q(
      \o_values[40] [2]), .QN());
   DFF_X1 \o_values_reg[40][1]  (.D(o_values[1]), .CK(n_0_127), .Q(
      \o_values[40] [1]), .QN());
   DFF_X1 \o_values_reg[40][0]  (.D(o_values[0]), .CK(n_0_127), .Q(
      \o_values[40] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[39]_reg  (.CK(clk), .E(n_0_44), .SE(1'b0), 
      .GCK(n_0_128));
   DFF_X1 \o_values_reg[39][15]  (.D(o_values[15]), .CK(n_0_128), .Q(
      \o_values[39] [15]), .QN());
   DFF_X1 \o_values_reg[39][14]  (.D(o_values[14]), .CK(n_0_128), .Q(
      \o_values[39] [14]), .QN());
   DFF_X1 \o_values_reg[39][13]  (.D(o_values[13]), .CK(n_0_128), .Q(
      \o_values[39] [13]), .QN());
   DFF_X1 \o_values_reg[39][12]  (.D(o_values[12]), .CK(n_0_128), .Q(
      \o_values[39] [12]), .QN());
   DFF_X1 \o_values_reg[39][11]  (.D(o_values[11]), .CK(n_0_128), .Q(
      \o_values[39] [11]), .QN());
   DFF_X1 \o_values_reg[39][10]  (.D(o_values[10]), .CK(n_0_128), .Q(
      \o_values[39] [10]), .QN());
   DFF_X1 \o_values_reg[39][9]  (.D(o_values[9]), .CK(n_0_128), .Q(
      \o_values[39] [9]), .QN());
   DFF_X1 \o_values_reg[39][8]  (.D(o_values[8]), .CK(n_0_128), .Q(
      \o_values[39] [8]), .QN());
   DFF_X1 \o_values_reg[39][7]  (.D(o_values[7]), .CK(n_0_128), .Q(
      \o_values[39] [7]), .QN());
   DFF_X1 \o_values_reg[39][6]  (.D(o_values[6]), .CK(n_0_128), .Q(
      \o_values[39] [6]), .QN());
   DFF_X1 \o_values_reg[39][5]  (.D(o_values[5]), .CK(n_0_128), .Q(
      \o_values[39] [5]), .QN());
   DFF_X1 \o_values_reg[39][4]  (.D(o_values[4]), .CK(n_0_128), .Q(
      \o_values[39] [4]), .QN());
   DFF_X1 \o_values_reg[39][3]  (.D(o_values[3]), .CK(n_0_128), .Q(
      \o_values[39] [3]), .QN());
   DFF_X1 \o_values_reg[39][2]  (.D(o_values[2]), .CK(n_0_128), .Q(
      \o_values[39] [2]), .QN());
   DFF_X1 \o_values_reg[39][1]  (.D(o_values[1]), .CK(n_0_128), .Q(
      \o_values[39] [1]), .QN());
   DFF_X1 \o_values_reg[39][0]  (.D(o_values[0]), .CK(n_0_128), .Q(
      \o_values[39] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[38]_reg  (.CK(clk), .E(n_0_45), .SE(1'b0), 
      .GCK(n_0_129));
   DFF_X1 \o_values_reg[38][15]  (.D(o_values[15]), .CK(n_0_129), .Q(
      \o_values[38] [15]), .QN());
   DFF_X1 \o_values_reg[38][14]  (.D(o_values[14]), .CK(n_0_129), .Q(
      \o_values[38] [14]), .QN());
   DFF_X1 \o_values_reg[38][13]  (.D(o_values[13]), .CK(n_0_129), .Q(
      \o_values[38] [13]), .QN());
   DFF_X1 \o_values_reg[38][12]  (.D(o_values[12]), .CK(n_0_129), .Q(
      \o_values[38] [12]), .QN());
   DFF_X1 \o_values_reg[38][11]  (.D(o_values[11]), .CK(n_0_129), .Q(
      \o_values[38] [11]), .QN());
   DFF_X1 \o_values_reg[38][10]  (.D(o_values[10]), .CK(n_0_129), .Q(
      \o_values[38] [10]), .QN());
   DFF_X1 \o_values_reg[38][9]  (.D(o_values[9]), .CK(n_0_129), .Q(
      \o_values[38] [9]), .QN());
   DFF_X1 \o_values_reg[38][8]  (.D(o_values[8]), .CK(n_0_129), .Q(
      \o_values[38] [8]), .QN());
   DFF_X1 \o_values_reg[38][7]  (.D(o_values[7]), .CK(n_0_129), .Q(
      \o_values[38] [7]), .QN());
   DFF_X1 \o_values_reg[38][6]  (.D(o_values[6]), .CK(n_0_129), .Q(
      \o_values[38] [6]), .QN());
   DFF_X1 \o_values_reg[38][5]  (.D(o_values[5]), .CK(n_0_129), .Q(
      \o_values[38] [5]), .QN());
   DFF_X1 \o_values_reg[38][4]  (.D(o_values[4]), .CK(n_0_129), .Q(
      \o_values[38] [4]), .QN());
   DFF_X1 \o_values_reg[38][3]  (.D(o_values[3]), .CK(n_0_129), .Q(
      \o_values[38] [3]), .QN());
   DFF_X1 \o_values_reg[38][2]  (.D(o_values[2]), .CK(n_0_129), .Q(
      \o_values[38] [2]), .QN());
   DFF_X1 \o_values_reg[38][1]  (.D(o_values[1]), .CK(n_0_129), .Q(
      \o_values[38] [1]), .QN());
   DFF_X1 \o_values_reg[38][0]  (.D(o_values[0]), .CK(n_0_129), .Q(
      \o_values[38] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[37]_reg  (.CK(clk), .E(n_0_46), .SE(1'b0), 
      .GCK(n_0_130));
   DFF_X1 \o_values_reg[37][15]  (.D(o_values[15]), .CK(n_0_130), .Q(
      \o_values[37] [15]), .QN());
   DFF_X1 \o_values_reg[37][14]  (.D(o_values[14]), .CK(n_0_130), .Q(
      \o_values[37] [14]), .QN());
   DFF_X1 \o_values_reg[37][13]  (.D(o_values[13]), .CK(n_0_130), .Q(
      \o_values[37] [13]), .QN());
   DFF_X1 \o_values_reg[37][12]  (.D(o_values[12]), .CK(n_0_130), .Q(
      \o_values[37] [12]), .QN());
   DFF_X1 \o_values_reg[37][11]  (.D(o_values[11]), .CK(n_0_130), .Q(
      \o_values[37] [11]), .QN());
   DFF_X1 \o_values_reg[37][10]  (.D(o_values[10]), .CK(n_0_130), .Q(
      \o_values[37] [10]), .QN());
   DFF_X1 \o_values_reg[37][9]  (.D(o_values[9]), .CK(n_0_130), .Q(
      \o_values[37] [9]), .QN());
   DFF_X1 \o_values_reg[37][8]  (.D(o_values[8]), .CK(n_0_130), .Q(
      \o_values[37] [8]), .QN());
   DFF_X1 \o_values_reg[37][7]  (.D(o_values[7]), .CK(n_0_130), .Q(
      \o_values[37] [7]), .QN());
   DFF_X1 \o_values_reg[37][6]  (.D(o_values[6]), .CK(n_0_130), .Q(
      \o_values[37] [6]), .QN());
   DFF_X1 \o_values_reg[37][5]  (.D(o_values[5]), .CK(n_0_130), .Q(
      \o_values[37] [5]), .QN());
   DFF_X1 \o_values_reg[37][4]  (.D(o_values[4]), .CK(n_0_130), .Q(
      \o_values[37] [4]), .QN());
   DFF_X1 \o_values_reg[37][3]  (.D(o_values[3]), .CK(n_0_130), .Q(
      \o_values[37] [3]), .QN());
   DFF_X1 \o_values_reg[37][2]  (.D(o_values[2]), .CK(n_0_130), .Q(
      \o_values[37] [2]), .QN());
   DFF_X1 \o_values_reg[37][1]  (.D(o_values[1]), .CK(n_0_130), .Q(
      \o_values[37] [1]), .QN());
   DFF_X1 \o_values_reg[37][0]  (.D(o_values[0]), .CK(n_0_130), .Q(
      \o_values[37] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[36]_reg  (.CK(clk), .E(n_0_47), .SE(1'b0), 
      .GCK(n_0_131));
   DFF_X1 \o_values_reg[36][15]  (.D(o_values[15]), .CK(n_0_131), .Q(
      \o_values[36] [15]), .QN());
   DFF_X1 \o_values_reg[36][14]  (.D(o_values[14]), .CK(n_0_131), .Q(
      \o_values[36] [14]), .QN());
   DFF_X1 \o_values_reg[36][13]  (.D(o_values[13]), .CK(n_0_131), .Q(
      \o_values[36] [13]), .QN());
   DFF_X1 \o_values_reg[36][12]  (.D(o_values[12]), .CK(n_0_131), .Q(
      \o_values[36] [12]), .QN());
   DFF_X1 \o_values_reg[36][11]  (.D(o_values[11]), .CK(n_0_131), .Q(
      \o_values[36] [11]), .QN());
   DFF_X1 \o_values_reg[36][10]  (.D(o_values[10]), .CK(n_0_131), .Q(
      \o_values[36] [10]), .QN());
   DFF_X1 \o_values_reg[36][9]  (.D(o_values[9]), .CK(n_0_131), .Q(
      \o_values[36] [9]), .QN());
   DFF_X1 \o_values_reg[36][8]  (.D(o_values[8]), .CK(n_0_131), .Q(
      \o_values[36] [8]), .QN());
   DFF_X1 \o_values_reg[36][7]  (.D(o_values[7]), .CK(n_0_131), .Q(
      \o_values[36] [7]), .QN());
   DFF_X1 \o_values_reg[36][6]  (.D(o_values[6]), .CK(n_0_131), .Q(
      \o_values[36] [6]), .QN());
   DFF_X1 \o_values_reg[36][5]  (.D(o_values[5]), .CK(n_0_131), .Q(
      \o_values[36] [5]), .QN());
   DFF_X1 \o_values_reg[36][4]  (.D(o_values[4]), .CK(n_0_131), .Q(
      \o_values[36] [4]), .QN());
   DFF_X1 \o_values_reg[36][3]  (.D(o_values[3]), .CK(n_0_131), .Q(
      \o_values[36] [3]), .QN());
   DFF_X1 \o_values_reg[36][2]  (.D(o_values[2]), .CK(n_0_131), .Q(
      \o_values[36] [2]), .QN());
   DFF_X1 \o_values_reg[36][1]  (.D(o_values[1]), .CK(n_0_131), .Q(
      \o_values[36] [1]), .QN());
   DFF_X1 \o_values_reg[36][0]  (.D(o_values[0]), .CK(n_0_131), .Q(
      \o_values[36] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[35]_reg  (.CK(clk), .E(n_0_48), .SE(1'b0), 
      .GCK(n_0_132));
   DFF_X1 \o_values_reg[35][15]  (.D(o_values[15]), .CK(n_0_132), .Q(
      \o_values[35] [15]), .QN());
   DFF_X1 \o_values_reg[35][14]  (.D(o_values[14]), .CK(n_0_132), .Q(
      \o_values[35] [14]), .QN());
   DFF_X1 \o_values_reg[35][13]  (.D(o_values[13]), .CK(n_0_132), .Q(
      \o_values[35] [13]), .QN());
   DFF_X1 \o_values_reg[35][12]  (.D(o_values[12]), .CK(n_0_132), .Q(
      \o_values[35] [12]), .QN());
   DFF_X1 \o_values_reg[35][11]  (.D(o_values[11]), .CK(n_0_132), .Q(
      \o_values[35] [11]), .QN());
   DFF_X1 \o_values_reg[35][10]  (.D(o_values[10]), .CK(n_0_132), .Q(
      \o_values[35] [10]), .QN());
   DFF_X1 \o_values_reg[35][9]  (.D(o_values[9]), .CK(n_0_132), .Q(
      \o_values[35] [9]), .QN());
   DFF_X1 \o_values_reg[35][8]  (.D(o_values[8]), .CK(n_0_132), .Q(
      \o_values[35] [8]), .QN());
   DFF_X1 \o_values_reg[35][7]  (.D(o_values[7]), .CK(n_0_132), .Q(
      \o_values[35] [7]), .QN());
   DFF_X1 \o_values_reg[35][6]  (.D(o_values[6]), .CK(n_0_132), .Q(
      \o_values[35] [6]), .QN());
   DFF_X1 \o_values_reg[35][5]  (.D(o_values[5]), .CK(n_0_132), .Q(
      \o_values[35] [5]), .QN());
   DFF_X1 \o_values_reg[35][4]  (.D(o_values[4]), .CK(n_0_132), .Q(
      \o_values[35] [4]), .QN());
   DFF_X1 \o_values_reg[35][3]  (.D(o_values[3]), .CK(n_0_132), .Q(
      \o_values[35] [3]), .QN());
   DFF_X1 \o_values_reg[35][2]  (.D(o_values[2]), .CK(n_0_132), .Q(
      \o_values[35] [2]), .QN());
   DFF_X1 \o_values_reg[35][1]  (.D(o_values[1]), .CK(n_0_132), .Q(
      \o_values[35] [1]), .QN());
   DFF_X1 \o_values_reg[35][0]  (.D(o_values[0]), .CK(n_0_132), .Q(
      \o_values[35] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[34]_reg  (.CK(clk), .E(n_0_49), .SE(1'b0), 
      .GCK(n_0_133));
   DFF_X1 \o_values_reg[34][15]  (.D(o_values[15]), .CK(n_0_133), .Q(
      \o_values[34] [15]), .QN());
   DFF_X1 \o_values_reg[34][14]  (.D(o_values[14]), .CK(n_0_133), .Q(
      \o_values[34] [14]), .QN());
   DFF_X1 \o_values_reg[34][13]  (.D(o_values[13]), .CK(n_0_133), .Q(
      \o_values[34] [13]), .QN());
   DFF_X1 \o_values_reg[34][12]  (.D(o_values[12]), .CK(n_0_133), .Q(
      \o_values[34] [12]), .QN());
   DFF_X1 \o_values_reg[34][11]  (.D(o_values[11]), .CK(n_0_133), .Q(
      \o_values[34] [11]), .QN());
   DFF_X1 \o_values_reg[34][10]  (.D(o_values[10]), .CK(n_0_133), .Q(
      \o_values[34] [10]), .QN());
   DFF_X1 \o_values_reg[34][9]  (.D(o_values[9]), .CK(n_0_133), .Q(
      \o_values[34] [9]), .QN());
   DFF_X1 \o_values_reg[34][8]  (.D(o_values[8]), .CK(n_0_133), .Q(
      \o_values[34] [8]), .QN());
   DFF_X1 \o_values_reg[34][7]  (.D(o_values[7]), .CK(n_0_133), .Q(
      \o_values[34] [7]), .QN());
   DFF_X1 \o_values_reg[34][6]  (.D(o_values[6]), .CK(n_0_133), .Q(
      \o_values[34] [6]), .QN());
   DFF_X1 \o_values_reg[34][5]  (.D(o_values[5]), .CK(n_0_133), .Q(
      \o_values[34] [5]), .QN());
   DFF_X1 \o_values_reg[34][4]  (.D(o_values[4]), .CK(n_0_133), .Q(
      \o_values[34] [4]), .QN());
   DFF_X1 \o_values_reg[34][3]  (.D(o_values[3]), .CK(n_0_133), .Q(
      \o_values[34] [3]), .QN());
   DFF_X1 \o_values_reg[34][2]  (.D(o_values[2]), .CK(n_0_133), .Q(
      \o_values[34] [2]), .QN());
   DFF_X1 \o_values_reg[34][1]  (.D(o_values[1]), .CK(n_0_133), .Q(
      \o_values[34] [1]), .QN());
   DFF_X1 \o_values_reg[34][0]  (.D(o_values[0]), .CK(n_0_133), .Q(
      \o_values[34] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[33]_reg  (.CK(clk), .E(n_0_50), .SE(1'b0), 
      .GCK(n_0_134));
   DFF_X1 \o_values_reg[33][15]  (.D(o_values[15]), .CK(n_0_134), .Q(
      \o_values[33] [15]), .QN());
   DFF_X1 \o_values_reg[33][14]  (.D(o_values[14]), .CK(n_0_134), .Q(
      \o_values[33] [14]), .QN());
   DFF_X1 \o_values_reg[33][13]  (.D(o_values[13]), .CK(n_0_134), .Q(
      \o_values[33] [13]), .QN());
   DFF_X1 \o_values_reg[33][12]  (.D(o_values[12]), .CK(n_0_134), .Q(
      \o_values[33] [12]), .QN());
   DFF_X1 \o_values_reg[33][11]  (.D(o_values[11]), .CK(n_0_134), .Q(
      \o_values[33] [11]), .QN());
   DFF_X1 \o_values_reg[33][10]  (.D(o_values[10]), .CK(n_0_134), .Q(
      \o_values[33] [10]), .QN());
   DFF_X1 \o_values_reg[33][9]  (.D(o_values[9]), .CK(n_0_134), .Q(
      \o_values[33] [9]), .QN());
   DFF_X1 \o_values_reg[33][8]  (.D(o_values[8]), .CK(n_0_134), .Q(
      \o_values[33] [8]), .QN());
   DFF_X1 \o_values_reg[33][7]  (.D(o_values[7]), .CK(n_0_134), .Q(
      \o_values[33] [7]), .QN());
   DFF_X1 \o_values_reg[33][6]  (.D(o_values[6]), .CK(n_0_134), .Q(
      \o_values[33] [6]), .QN());
   DFF_X1 \o_values_reg[33][5]  (.D(o_values[5]), .CK(n_0_134), .Q(
      \o_values[33] [5]), .QN());
   DFF_X1 \o_values_reg[33][4]  (.D(o_values[4]), .CK(n_0_134), .Q(
      \o_values[33] [4]), .QN());
   DFF_X1 \o_values_reg[33][3]  (.D(o_values[3]), .CK(n_0_134), .Q(
      \o_values[33] [3]), .QN());
   DFF_X1 \o_values_reg[33][2]  (.D(o_values[2]), .CK(n_0_134), .Q(
      \o_values[33] [2]), .QN());
   DFF_X1 \o_values_reg[33][1]  (.D(o_values[1]), .CK(n_0_134), .Q(
      \o_values[33] [1]), .QN());
   DFF_X1 \o_values_reg[33][0]  (.D(o_values[0]), .CK(n_0_134), .Q(
      \o_values[33] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[32]_reg  (.CK(clk), .E(n_0_51), .SE(1'b0), 
      .GCK(n_0_135));
   DFF_X1 \o_values_reg[32][15]  (.D(o_values[15]), .CK(n_0_135), .Q(
      \o_values[32] [15]), .QN());
   DFF_X1 \o_values_reg[32][14]  (.D(o_values[14]), .CK(n_0_135), .Q(
      \o_values[32] [14]), .QN());
   DFF_X1 \o_values_reg[32][13]  (.D(o_values[13]), .CK(n_0_135), .Q(
      \o_values[32] [13]), .QN());
   DFF_X1 \o_values_reg[32][12]  (.D(o_values[12]), .CK(n_0_135), .Q(
      \o_values[32] [12]), .QN());
   DFF_X1 \o_values_reg[32][11]  (.D(o_values[11]), .CK(n_0_135), .Q(
      \o_values[32] [11]), .QN());
   DFF_X1 \o_values_reg[32][10]  (.D(o_values[10]), .CK(n_0_135), .Q(
      \o_values[32] [10]), .QN());
   DFF_X1 \o_values_reg[32][9]  (.D(o_values[9]), .CK(n_0_135), .Q(
      \o_values[32] [9]), .QN());
   DFF_X1 \o_values_reg[32][8]  (.D(o_values[8]), .CK(n_0_135), .Q(
      \o_values[32] [8]), .QN());
   DFF_X1 \o_values_reg[32][7]  (.D(o_values[7]), .CK(n_0_135), .Q(
      \o_values[32] [7]), .QN());
   DFF_X1 \o_values_reg[32][6]  (.D(o_values[6]), .CK(n_0_135), .Q(
      \o_values[32] [6]), .QN());
   DFF_X1 \o_values_reg[32][5]  (.D(o_values[5]), .CK(n_0_135), .Q(
      \o_values[32] [5]), .QN());
   DFF_X1 \o_values_reg[32][4]  (.D(o_values[4]), .CK(n_0_135), .Q(
      \o_values[32] [4]), .QN());
   DFF_X1 \o_values_reg[32][3]  (.D(o_values[3]), .CK(n_0_135), .Q(
      \o_values[32] [3]), .QN());
   DFF_X1 \o_values_reg[32][2]  (.D(o_values[2]), .CK(n_0_135), .Q(
      \o_values[32] [2]), .QN());
   DFF_X1 \o_values_reg[32][1]  (.D(o_values[1]), .CK(n_0_135), .Q(
      \o_values[32] [1]), .QN());
   DFF_X1 \o_values_reg[32][0]  (.D(o_values[0]), .CK(n_0_135), .Q(
      \o_values[32] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[31]_reg  (.CK(clk), .E(n_0_52), .SE(1'b0), 
      .GCK(n_0_136));
   DFF_X1 \o_values_reg[31][15]  (.D(o_values[15]), .CK(n_0_136), .Q(
      \o_values[31] [15]), .QN());
   DFF_X1 \o_values_reg[31][14]  (.D(o_values[14]), .CK(n_0_136), .Q(
      \o_values[31] [14]), .QN());
   DFF_X1 \o_values_reg[31][13]  (.D(o_values[13]), .CK(n_0_136), .Q(
      \o_values[31] [13]), .QN());
   DFF_X1 \o_values_reg[31][12]  (.D(o_values[12]), .CK(n_0_136), .Q(
      \o_values[31] [12]), .QN());
   DFF_X1 \o_values_reg[31][11]  (.D(o_values[11]), .CK(n_0_136), .Q(
      \o_values[31] [11]), .QN());
   DFF_X1 \o_values_reg[31][10]  (.D(o_values[10]), .CK(n_0_136), .Q(
      \o_values[31] [10]), .QN());
   DFF_X1 \o_values_reg[31][9]  (.D(o_values[9]), .CK(n_0_136), .Q(
      \o_values[31] [9]), .QN());
   DFF_X1 \o_values_reg[31][8]  (.D(o_values[8]), .CK(n_0_136), .Q(
      \o_values[31] [8]), .QN());
   DFF_X1 \o_values_reg[31][7]  (.D(o_values[7]), .CK(n_0_136), .Q(
      \o_values[31] [7]), .QN());
   DFF_X1 \o_values_reg[31][6]  (.D(o_values[6]), .CK(n_0_136), .Q(
      \o_values[31] [6]), .QN());
   DFF_X1 \o_values_reg[31][5]  (.D(o_values[5]), .CK(n_0_136), .Q(
      \o_values[31] [5]), .QN());
   DFF_X1 \o_values_reg[31][4]  (.D(o_values[4]), .CK(n_0_136), .Q(
      \o_values[31] [4]), .QN());
   DFF_X1 \o_values_reg[31][3]  (.D(o_values[3]), .CK(n_0_136), .Q(
      \o_values[31] [3]), .QN());
   DFF_X1 \o_values_reg[31][2]  (.D(o_values[2]), .CK(n_0_136), .Q(
      \o_values[31] [2]), .QN());
   DFF_X1 \o_values_reg[31][1]  (.D(o_values[1]), .CK(n_0_136), .Q(
      \o_values[31] [1]), .QN());
   DFF_X1 \o_values_reg[31][0]  (.D(o_values[0]), .CK(n_0_136), .Q(
      \o_values[31] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[30]_reg  (.CK(clk), .E(n_0_53), .SE(1'b0), 
      .GCK(n_0_137));
   DFF_X1 \o_values_reg[30][15]  (.D(o_values[15]), .CK(n_0_137), .Q(
      \o_values[30] [15]), .QN());
   DFF_X1 \o_values_reg[30][14]  (.D(o_values[14]), .CK(n_0_137), .Q(
      \o_values[30] [14]), .QN());
   DFF_X1 \o_values_reg[30][13]  (.D(o_values[13]), .CK(n_0_137), .Q(
      \o_values[30] [13]), .QN());
   DFF_X1 \o_values_reg[30][12]  (.D(o_values[12]), .CK(n_0_137), .Q(
      \o_values[30] [12]), .QN());
   DFF_X1 \o_values_reg[30][11]  (.D(o_values[11]), .CK(n_0_137), .Q(
      \o_values[30] [11]), .QN());
   DFF_X1 \o_values_reg[30][10]  (.D(o_values[10]), .CK(n_0_137), .Q(
      \o_values[30] [10]), .QN());
   DFF_X1 \o_values_reg[30][9]  (.D(o_values[9]), .CK(n_0_137), .Q(
      \o_values[30] [9]), .QN());
   DFF_X1 \o_values_reg[30][8]  (.D(o_values[8]), .CK(n_0_137), .Q(
      \o_values[30] [8]), .QN());
   DFF_X1 \o_values_reg[30][7]  (.D(o_values[7]), .CK(n_0_137), .Q(
      \o_values[30] [7]), .QN());
   DFF_X1 \o_values_reg[30][6]  (.D(o_values[6]), .CK(n_0_137), .Q(
      \o_values[30] [6]), .QN());
   DFF_X1 \o_values_reg[30][5]  (.D(o_values[5]), .CK(n_0_137), .Q(
      \o_values[30] [5]), .QN());
   DFF_X1 \o_values_reg[30][4]  (.D(o_values[4]), .CK(n_0_137), .Q(
      \o_values[30] [4]), .QN());
   DFF_X1 \o_values_reg[30][3]  (.D(o_values[3]), .CK(n_0_137), .Q(
      \o_values[30] [3]), .QN());
   DFF_X1 \o_values_reg[30][2]  (.D(o_values[2]), .CK(n_0_137), .Q(
      \o_values[30] [2]), .QN());
   DFF_X1 \o_values_reg[30][1]  (.D(o_values[1]), .CK(n_0_137), .Q(
      \o_values[30] [1]), .QN());
   DFF_X1 \o_values_reg[30][0]  (.D(o_values[0]), .CK(n_0_137), .Q(
      \o_values[30] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[29]_reg  (.CK(clk), .E(n_0_54), .SE(1'b0), 
      .GCK(n_0_138));
   DFF_X1 \o_values_reg[29][15]  (.D(o_values[15]), .CK(n_0_138), .Q(
      \o_values[29] [15]), .QN());
   DFF_X1 \o_values_reg[29][14]  (.D(o_values[14]), .CK(n_0_138), .Q(
      \o_values[29] [14]), .QN());
   DFF_X1 \o_values_reg[29][13]  (.D(o_values[13]), .CK(n_0_138), .Q(
      \o_values[29] [13]), .QN());
   DFF_X1 \o_values_reg[29][12]  (.D(o_values[12]), .CK(n_0_138), .Q(
      \o_values[29] [12]), .QN());
   DFF_X1 \o_values_reg[29][11]  (.D(o_values[11]), .CK(n_0_138), .Q(
      \o_values[29] [11]), .QN());
   DFF_X1 \o_values_reg[29][10]  (.D(o_values[10]), .CK(n_0_138), .Q(
      \o_values[29] [10]), .QN());
   DFF_X1 \o_values_reg[29][9]  (.D(o_values[9]), .CK(n_0_138), .Q(
      \o_values[29] [9]), .QN());
   DFF_X1 \o_values_reg[29][8]  (.D(o_values[8]), .CK(n_0_138), .Q(
      \o_values[29] [8]), .QN());
   DFF_X1 \o_values_reg[29][7]  (.D(o_values[7]), .CK(n_0_138), .Q(
      \o_values[29] [7]), .QN());
   DFF_X1 \o_values_reg[29][6]  (.D(o_values[6]), .CK(n_0_138), .Q(
      \o_values[29] [6]), .QN());
   DFF_X1 \o_values_reg[29][5]  (.D(o_values[5]), .CK(n_0_138), .Q(
      \o_values[29] [5]), .QN());
   DFF_X1 \o_values_reg[29][4]  (.D(o_values[4]), .CK(n_0_138), .Q(
      \o_values[29] [4]), .QN());
   DFF_X1 \o_values_reg[29][3]  (.D(o_values[3]), .CK(n_0_138), .Q(
      \o_values[29] [3]), .QN());
   DFF_X1 \o_values_reg[29][2]  (.D(o_values[2]), .CK(n_0_138), .Q(
      \o_values[29] [2]), .QN());
   DFF_X1 \o_values_reg[29][1]  (.D(o_values[1]), .CK(n_0_138), .Q(
      \o_values[29] [1]), .QN());
   DFF_X1 \o_values_reg[29][0]  (.D(o_values[0]), .CK(n_0_138), .Q(
      \o_values[29] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[28]_reg  (.CK(clk), .E(n_0_55), .SE(1'b0), 
      .GCK(n_0_139));
   DFF_X1 \o_values_reg[28][15]  (.D(o_values[15]), .CK(n_0_139), .Q(
      \o_values[28] [15]), .QN());
   DFF_X1 \o_values_reg[28][14]  (.D(o_values[14]), .CK(n_0_139), .Q(
      \o_values[28] [14]), .QN());
   DFF_X1 \o_values_reg[28][13]  (.D(o_values[13]), .CK(n_0_139), .Q(
      \o_values[28] [13]), .QN());
   DFF_X1 \o_values_reg[28][12]  (.D(o_values[12]), .CK(n_0_139), .Q(
      \o_values[28] [12]), .QN());
   DFF_X1 \o_values_reg[28][11]  (.D(o_values[11]), .CK(n_0_139), .Q(
      \o_values[28] [11]), .QN());
   DFF_X1 \o_values_reg[28][10]  (.D(o_values[10]), .CK(n_0_139), .Q(
      \o_values[28] [10]), .QN());
   DFF_X1 \o_values_reg[28][9]  (.D(o_values[9]), .CK(n_0_139), .Q(
      \o_values[28] [9]), .QN());
   DFF_X1 \o_values_reg[28][8]  (.D(o_values[8]), .CK(n_0_139), .Q(
      \o_values[28] [8]), .QN());
   DFF_X1 \o_values_reg[28][7]  (.D(o_values[7]), .CK(n_0_139), .Q(
      \o_values[28] [7]), .QN());
   DFF_X1 \o_values_reg[28][6]  (.D(o_values[6]), .CK(n_0_139), .Q(
      \o_values[28] [6]), .QN());
   DFF_X1 \o_values_reg[28][5]  (.D(o_values[5]), .CK(n_0_139), .Q(
      \o_values[28] [5]), .QN());
   DFF_X1 \o_values_reg[28][4]  (.D(o_values[4]), .CK(n_0_139), .Q(
      \o_values[28] [4]), .QN());
   DFF_X1 \o_values_reg[28][3]  (.D(o_values[3]), .CK(n_0_139), .Q(
      \o_values[28] [3]), .QN());
   DFF_X1 \o_values_reg[28][2]  (.D(o_values[2]), .CK(n_0_139), .Q(
      \o_values[28] [2]), .QN());
   DFF_X1 \o_values_reg[28][1]  (.D(o_values[1]), .CK(n_0_139), .Q(
      \o_values[28] [1]), .QN());
   DFF_X1 \o_values_reg[28][0]  (.D(o_values[0]), .CK(n_0_139), .Q(
      \o_values[28] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[27]_reg  (.CK(clk), .E(n_0_56), .SE(1'b0), 
      .GCK(n_0_140));
   DFF_X1 \o_values_reg[27][15]  (.D(o_values[15]), .CK(n_0_140), .Q(
      \o_values[27] [15]), .QN());
   DFF_X1 \o_values_reg[27][14]  (.D(o_values[14]), .CK(n_0_140), .Q(
      \o_values[27] [14]), .QN());
   DFF_X1 \o_values_reg[27][13]  (.D(o_values[13]), .CK(n_0_140), .Q(
      \o_values[27] [13]), .QN());
   DFF_X1 \o_values_reg[27][12]  (.D(o_values[12]), .CK(n_0_140), .Q(
      \o_values[27] [12]), .QN());
   DFF_X1 \o_values_reg[27][11]  (.D(o_values[11]), .CK(n_0_140), .Q(
      \o_values[27] [11]), .QN());
   DFF_X1 \o_values_reg[27][10]  (.D(o_values[10]), .CK(n_0_140), .Q(
      \o_values[27] [10]), .QN());
   DFF_X1 \o_values_reg[27][9]  (.D(o_values[9]), .CK(n_0_140), .Q(
      \o_values[27] [9]), .QN());
   DFF_X1 \o_values_reg[27][8]  (.D(o_values[8]), .CK(n_0_140), .Q(
      \o_values[27] [8]), .QN());
   DFF_X1 \o_values_reg[27][7]  (.D(o_values[7]), .CK(n_0_140), .Q(
      \o_values[27] [7]), .QN());
   DFF_X1 \o_values_reg[27][6]  (.D(o_values[6]), .CK(n_0_140), .Q(
      \o_values[27] [6]), .QN());
   DFF_X1 \o_values_reg[27][5]  (.D(o_values[5]), .CK(n_0_140), .Q(
      \o_values[27] [5]), .QN());
   DFF_X1 \o_values_reg[27][4]  (.D(o_values[4]), .CK(n_0_140), .Q(
      \o_values[27] [4]), .QN());
   DFF_X1 \o_values_reg[27][3]  (.D(o_values[3]), .CK(n_0_140), .Q(
      \o_values[27] [3]), .QN());
   DFF_X1 \o_values_reg[27][2]  (.D(o_values[2]), .CK(n_0_140), .Q(
      \o_values[27] [2]), .QN());
   DFF_X1 \o_values_reg[27][1]  (.D(o_values[1]), .CK(n_0_140), .Q(
      \o_values[27] [1]), .QN());
   DFF_X1 \o_values_reg[27][0]  (.D(o_values[0]), .CK(n_0_140), .Q(
      \o_values[27] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[26]_reg  (.CK(clk), .E(n_0_57), .SE(1'b0), 
      .GCK(n_0_141));
   DFF_X1 \o_values_reg[26][15]  (.D(o_values[15]), .CK(n_0_141), .Q(
      \o_values[26] [15]), .QN());
   DFF_X1 \o_values_reg[26][14]  (.D(o_values[14]), .CK(n_0_141), .Q(
      \o_values[26] [14]), .QN());
   DFF_X1 \o_values_reg[26][13]  (.D(o_values[13]), .CK(n_0_141), .Q(
      \o_values[26] [13]), .QN());
   DFF_X1 \o_values_reg[26][12]  (.D(o_values[12]), .CK(n_0_141), .Q(
      \o_values[26] [12]), .QN());
   DFF_X1 \o_values_reg[26][11]  (.D(o_values[11]), .CK(n_0_141), .Q(
      \o_values[26] [11]), .QN());
   DFF_X1 \o_values_reg[26][10]  (.D(o_values[10]), .CK(n_0_141), .Q(
      \o_values[26] [10]), .QN());
   DFF_X1 \o_values_reg[26][9]  (.D(o_values[9]), .CK(n_0_141), .Q(
      \o_values[26] [9]), .QN());
   DFF_X1 \o_values_reg[26][8]  (.D(o_values[8]), .CK(n_0_141), .Q(
      \o_values[26] [8]), .QN());
   DFF_X1 \o_values_reg[26][7]  (.D(o_values[7]), .CK(n_0_141), .Q(
      \o_values[26] [7]), .QN());
   DFF_X1 \o_values_reg[26][6]  (.D(o_values[6]), .CK(n_0_141), .Q(
      \o_values[26] [6]), .QN());
   DFF_X1 \o_values_reg[26][5]  (.D(o_values[5]), .CK(n_0_141), .Q(
      \o_values[26] [5]), .QN());
   DFF_X1 \o_values_reg[26][4]  (.D(o_values[4]), .CK(n_0_141), .Q(
      \o_values[26] [4]), .QN());
   DFF_X1 \o_values_reg[26][3]  (.D(o_values[3]), .CK(n_0_141), .Q(
      \o_values[26] [3]), .QN());
   DFF_X1 \o_values_reg[26][2]  (.D(o_values[2]), .CK(n_0_141), .Q(
      \o_values[26] [2]), .QN());
   DFF_X1 \o_values_reg[26][1]  (.D(o_values[1]), .CK(n_0_141), .Q(
      \o_values[26] [1]), .QN());
   DFF_X1 \o_values_reg[26][0]  (.D(o_values[0]), .CK(n_0_141), .Q(
      \o_values[26] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[25]_reg  (.CK(clk), .E(n_0_58), .SE(1'b0), 
      .GCK(n_0_142));
   DFF_X1 \o_values_reg[25][15]  (.D(o_values[15]), .CK(n_0_142), .Q(
      \o_values[25] [15]), .QN());
   DFF_X1 \o_values_reg[25][14]  (.D(o_values[14]), .CK(n_0_142), .Q(
      \o_values[25] [14]), .QN());
   DFF_X1 \o_values_reg[25][13]  (.D(o_values[13]), .CK(n_0_142), .Q(
      \o_values[25] [13]), .QN());
   DFF_X1 \o_values_reg[25][12]  (.D(o_values[12]), .CK(n_0_142), .Q(
      \o_values[25] [12]), .QN());
   DFF_X1 \o_values_reg[25][11]  (.D(o_values[11]), .CK(n_0_142), .Q(
      \o_values[25] [11]), .QN());
   DFF_X1 \o_values_reg[25][10]  (.D(o_values[10]), .CK(n_0_142), .Q(
      \o_values[25] [10]), .QN());
   DFF_X1 \o_values_reg[25][9]  (.D(o_values[9]), .CK(n_0_142), .Q(
      \o_values[25] [9]), .QN());
   DFF_X1 \o_values_reg[25][8]  (.D(o_values[8]), .CK(n_0_142), .Q(
      \o_values[25] [8]), .QN());
   DFF_X1 \o_values_reg[25][7]  (.D(o_values[7]), .CK(n_0_142), .Q(
      \o_values[25] [7]), .QN());
   DFF_X1 \o_values_reg[25][6]  (.D(o_values[6]), .CK(n_0_142), .Q(
      \o_values[25] [6]), .QN());
   DFF_X1 \o_values_reg[25][5]  (.D(o_values[5]), .CK(n_0_142), .Q(
      \o_values[25] [5]), .QN());
   DFF_X1 \o_values_reg[25][4]  (.D(o_values[4]), .CK(n_0_142), .Q(
      \o_values[25] [4]), .QN());
   DFF_X1 \o_values_reg[25][3]  (.D(o_values[3]), .CK(n_0_142), .Q(
      \o_values[25] [3]), .QN());
   DFF_X1 \o_values_reg[25][2]  (.D(o_values[2]), .CK(n_0_142), .Q(
      \o_values[25] [2]), .QN());
   DFF_X1 \o_values_reg[25][1]  (.D(o_values[1]), .CK(n_0_142), .Q(
      \o_values[25] [1]), .QN());
   DFF_X1 \o_values_reg[25][0]  (.D(o_values[0]), .CK(n_0_142), .Q(
      \o_values[25] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[24]_reg  (.CK(clk), .E(n_0_59), .SE(1'b0), 
      .GCK(n_0_143));
   DFF_X1 \o_values_reg[24][15]  (.D(o_values[15]), .CK(n_0_143), .Q(
      \o_values[24] [15]), .QN());
   DFF_X1 \o_values_reg[24][14]  (.D(o_values[14]), .CK(n_0_143), .Q(
      \o_values[24] [14]), .QN());
   DFF_X1 \o_values_reg[24][13]  (.D(o_values[13]), .CK(n_0_143), .Q(
      \o_values[24] [13]), .QN());
   DFF_X1 \o_values_reg[24][12]  (.D(o_values[12]), .CK(n_0_143), .Q(
      \o_values[24] [12]), .QN());
   DFF_X1 \o_values_reg[24][11]  (.D(o_values[11]), .CK(n_0_143), .Q(
      \o_values[24] [11]), .QN());
   DFF_X1 \o_values_reg[24][10]  (.D(o_values[10]), .CK(n_0_143), .Q(
      \o_values[24] [10]), .QN());
   DFF_X1 \o_values_reg[24][9]  (.D(o_values[9]), .CK(n_0_143), .Q(
      \o_values[24] [9]), .QN());
   DFF_X1 \o_values_reg[24][8]  (.D(o_values[8]), .CK(n_0_143), .Q(
      \o_values[24] [8]), .QN());
   DFF_X1 \o_values_reg[24][7]  (.D(o_values[7]), .CK(n_0_143), .Q(
      \o_values[24] [7]), .QN());
   DFF_X1 \o_values_reg[24][6]  (.D(o_values[6]), .CK(n_0_143), .Q(
      \o_values[24] [6]), .QN());
   DFF_X1 \o_values_reg[24][5]  (.D(o_values[5]), .CK(n_0_143), .Q(
      \o_values[24] [5]), .QN());
   DFF_X1 \o_values_reg[24][4]  (.D(o_values[4]), .CK(n_0_143), .Q(
      \o_values[24] [4]), .QN());
   DFF_X1 \o_values_reg[24][3]  (.D(o_values[3]), .CK(n_0_143), .Q(
      \o_values[24] [3]), .QN());
   DFF_X1 \o_values_reg[24][2]  (.D(o_values[2]), .CK(n_0_143), .Q(
      \o_values[24] [2]), .QN());
   DFF_X1 \o_values_reg[24][1]  (.D(o_values[1]), .CK(n_0_143), .Q(
      \o_values[24] [1]), .QN());
   DFF_X1 \o_values_reg[24][0]  (.D(o_values[0]), .CK(n_0_143), .Q(
      \o_values[24] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[23]_reg  (.CK(clk), .E(n_0_60), .SE(1'b0), 
      .GCK(n_0_144));
   DFF_X1 \o_values_reg[23][15]  (.D(o_values[15]), .CK(n_0_144), .Q(
      \o_values[23] [15]), .QN());
   DFF_X1 \o_values_reg[23][14]  (.D(o_values[14]), .CK(n_0_144), .Q(
      \o_values[23] [14]), .QN());
   DFF_X1 \o_values_reg[23][13]  (.D(o_values[13]), .CK(n_0_144), .Q(
      \o_values[23] [13]), .QN());
   DFF_X1 \o_values_reg[23][12]  (.D(o_values[12]), .CK(n_0_144), .Q(
      \o_values[23] [12]), .QN());
   DFF_X1 \o_values_reg[23][11]  (.D(o_values[11]), .CK(n_0_144), .Q(
      \o_values[23] [11]), .QN());
   DFF_X1 \o_values_reg[23][10]  (.D(o_values[10]), .CK(n_0_144), .Q(
      \o_values[23] [10]), .QN());
   DFF_X1 \o_values_reg[23][9]  (.D(o_values[9]), .CK(n_0_144), .Q(
      \o_values[23] [9]), .QN());
   DFF_X1 \o_values_reg[23][8]  (.D(o_values[8]), .CK(n_0_144), .Q(
      \o_values[23] [8]), .QN());
   DFF_X1 \o_values_reg[23][7]  (.D(o_values[7]), .CK(n_0_144), .Q(
      \o_values[23] [7]), .QN());
   DFF_X1 \o_values_reg[23][6]  (.D(o_values[6]), .CK(n_0_144), .Q(
      \o_values[23] [6]), .QN());
   DFF_X1 \o_values_reg[23][5]  (.D(o_values[5]), .CK(n_0_144), .Q(
      \o_values[23] [5]), .QN());
   DFF_X1 \o_values_reg[23][4]  (.D(o_values[4]), .CK(n_0_144), .Q(
      \o_values[23] [4]), .QN());
   DFF_X1 \o_values_reg[23][3]  (.D(o_values[3]), .CK(n_0_144), .Q(
      \o_values[23] [3]), .QN());
   DFF_X1 \o_values_reg[23][2]  (.D(o_values[2]), .CK(n_0_144), .Q(
      \o_values[23] [2]), .QN());
   DFF_X1 \o_values_reg[23][1]  (.D(o_values[1]), .CK(n_0_144), .Q(
      \o_values[23] [1]), .QN());
   DFF_X1 \o_values_reg[23][0]  (.D(o_values[0]), .CK(n_0_144), .Q(
      \o_values[23] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[22]_reg  (.CK(clk), .E(n_0_61), .SE(1'b0), 
      .GCK(n_0_145));
   DFF_X1 \o_values_reg[22][15]  (.D(o_values[15]), .CK(n_0_145), .Q(
      \o_values[22] [15]), .QN());
   DFF_X1 \o_values_reg[22][14]  (.D(o_values[14]), .CK(n_0_145), .Q(
      \o_values[22] [14]), .QN());
   DFF_X1 \o_values_reg[22][13]  (.D(o_values[13]), .CK(n_0_145), .Q(
      \o_values[22] [13]), .QN());
   DFF_X1 \o_values_reg[22][12]  (.D(o_values[12]), .CK(n_0_145), .Q(
      \o_values[22] [12]), .QN());
   DFF_X1 \o_values_reg[22][11]  (.D(o_values[11]), .CK(n_0_145), .Q(
      \o_values[22] [11]), .QN());
   DFF_X1 \o_values_reg[22][10]  (.D(o_values[10]), .CK(n_0_145), .Q(
      \o_values[22] [10]), .QN());
   DFF_X1 \o_values_reg[22][9]  (.D(o_values[9]), .CK(n_0_145), .Q(
      \o_values[22] [9]), .QN());
   DFF_X1 \o_values_reg[22][8]  (.D(o_values[8]), .CK(n_0_145), .Q(
      \o_values[22] [8]), .QN());
   DFF_X1 \o_values_reg[22][7]  (.D(o_values[7]), .CK(n_0_145), .Q(
      \o_values[22] [7]), .QN());
   DFF_X1 \o_values_reg[22][6]  (.D(o_values[6]), .CK(n_0_145), .Q(
      \o_values[22] [6]), .QN());
   DFF_X1 \o_values_reg[22][5]  (.D(o_values[5]), .CK(n_0_145), .Q(
      \o_values[22] [5]), .QN());
   DFF_X1 \o_values_reg[22][4]  (.D(o_values[4]), .CK(n_0_145), .Q(
      \o_values[22] [4]), .QN());
   DFF_X1 \o_values_reg[22][3]  (.D(o_values[3]), .CK(n_0_145), .Q(
      \o_values[22] [3]), .QN());
   DFF_X1 \o_values_reg[22][2]  (.D(o_values[2]), .CK(n_0_145), .Q(
      \o_values[22] [2]), .QN());
   DFF_X1 \o_values_reg[22][1]  (.D(o_values[1]), .CK(n_0_145), .Q(
      \o_values[22] [1]), .QN());
   DFF_X1 \o_values_reg[22][0]  (.D(o_values[0]), .CK(n_0_145), .Q(
      \o_values[22] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[21]_reg  (.CK(clk), .E(n_0_62), .SE(1'b0), 
      .GCK(n_0_146));
   DFF_X1 \o_values_reg[21][15]  (.D(o_values[15]), .CK(n_0_146), .Q(
      \o_values[21] [15]), .QN());
   DFF_X1 \o_values_reg[21][14]  (.D(o_values[14]), .CK(n_0_146), .Q(
      \o_values[21] [14]), .QN());
   DFF_X1 \o_values_reg[21][13]  (.D(o_values[13]), .CK(n_0_146), .Q(
      \o_values[21] [13]), .QN());
   DFF_X1 \o_values_reg[21][12]  (.D(o_values[12]), .CK(n_0_146), .Q(
      \o_values[21] [12]), .QN());
   DFF_X1 \o_values_reg[21][11]  (.D(o_values[11]), .CK(n_0_146), .Q(
      \o_values[21] [11]), .QN());
   DFF_X1 \o_values_reg[21][10]  (.D(o_values[10]), .CK(n_0_146), .Q(
      \o_values[21] [10]), .QN());
   DFF_X1 \o_values_reg[21][9]  (.D(o_values[9]), .CK(n_0_146), .Q(
      \o_values[21] [9]), .QN());
   DFF_X1 \o_values_reg[21][8]  (.D(o_values[8]), .CK(n_0_146), .Q(
      \o_values[21] [8]), .QN());
   DFF_X1 \o_values_reg[21][7]  (.D(o_values[7]), .CK(n_0_146), .Q(
      \o_values[21] [7]), .QN());
   DFF_X1 \o_values_reg[21][6]  (.D(o_values[6]), .CK(n_0_146), .Q(
      \o_values[21] [6]), .QN());
   DFF_X1 \o_values_reg[21][5]  (.D(o_values[5]), .CK(n_0_146), .Q(
      \o_values[21] [5]), .QN());
   DFF_X1 \o_values_reg[21][4]  (.D(o_values[4]), .CK(n_0_146), .Q(
      \o_values[21] [4]), .QN());
   DFF_X1 \o_values_reg[21][3]  (.D(o_values[3]), .CK(n_0_146), .Q(
      \o_values[21] [3]), .QN());
   DFF_X1 \o_values_reg[21][2]  (.D(o_values[2]), .CK(n_0_146), .Q(
      \o_values[21] [2]), .QN());
   DFF_X1 \o_values_reg[21][1]  (.D(o_values[1]), .CK(n_0_146), .Q(
      \o_values[21] [1]), .QN());
   DFF_X1 \o_values_reg[21][0]  (.D(o_values[0]), .CK(n_0_146), .Q(
      \o_values[21] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[20]_reg  (.CK(clk), .E(n_0_63), .SE(1'b0), 
      .GCK(n_0_147));
   DFF_X1 \o_values_reg[20][15]  (.D(o_values[15]), .CK(n_0_147), .Q(
      \o_values[20] [15]), .QN());
   DFF_X1 \o_values_reg[20][14]  (.D(o_values[14]), .CK(n_0_147), .Q(
      \o_values[20] [14]), .QN());
   DFF_X1 \o_values_reg[20][13]  (.D(o_values[13]), .CK(n_0_147), .Q(
      \o_values[20] [13]), .QN());
   DFF_X1 \o_values_reg[20][12]  (.D(o_values[12]), .CK(n_0_147), .Q(
      \o_values[20] [12]), .QN());
   DFF_X1 \o_values_reg[20][11]  (.D(o_values[11]), .CK(n_0_147), .Q(
      \o_values[20] [11]), .QN());
   DFF_X1 \o_values_reg[20][10]  (.D(o_values[10]), .CK(n_0_147), .Q(
      \o_values[20] [10]), .QN());
   DFF_X1 \o_values_reg[20][9]  (.D(o_values[9]), .CK(n_0_147), .Q(
      \o_values[20] [9]), .QN());
   DFF_X1 \o_values_reg[20][8]  (.D(o_values[8]), .CK(n_0_147), .Q(
      \o_values[20] [8]), .QN());
   DFF_X1 \o_values_reg[20][7]  (.D(o_values[7]), .CK(n_0_147), .Q(
      \o_values[20] [7]), .QN());
   DFF_X1 \o_values_reg[20][6]  (.D(o_values[6]), .CK(n_0_147), .Q(
      \o_values[20] [6]), .QN());
   DFF_X1 \o_values_reg[20][5]  (.D(o_values[5]), .CK(n_0_147), .Q(
      \o_values[20] [5]), .QN());
   DFF_X1 \o_values_reg[20][4]  (.D(o_values[4]), .CK(n_0_147), .Q(
      \o_values[20] [4]), .QN());
   DFF_X1 \o_values_reg[20][3]  (.D(o_values[3]), .CK(n_0_147), .Q(
      \o_values[20] [3]), .QN());
   DFF_X1 \o_values_reg[20][2]  (.D(o_values[2]), .CK(n_0_147), .Q(
      \o_values[20] [2]), .QN());
   DFF_X1 \o_values_reg[20][1]  (.D(o_values[1]), .CK(n_0_147), .Q(
      \o_values[20] [1]), .QN());
   DFF_X1 \o_values_reg[20][0]  (.D(o_values[0]), .CK(n_0_147), .Q(
      \o_values[20] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[19]_reg  (.CK(clk), .E(n_0_64), .SE(1'b0), 
      .GCK(n_0_148));
   DFF_X1 \o_values_reg[19][15]  (.D(o_values[15]), .CK(n_0_148), .Q(
      \o_values[19] [15]), .QN());
   DFF_X1 \o_values_reg[19][14]  (.D(o_values[14]), .CK(n_0_148), .Q(
      \o_values[19] [14]), .QN());
   DFF_X1 \o_values_reg[19][13]  (.D(o_values[13]), .CK(n_0_148), .Q(
      \o_values[19] [13]), .QN());
   DFF_X1 \o_values_reg[19][12]  (.D(o_values[12]), .CK(n_0_148), .Q(
      \o_values[19] [12]), .QN());
   DFF_X1 \o_values_reg[19][11]  (.D(o_values[11]), .CK(n_0_148), .Q(
      \o_values[19] [11]), .QN());
   DFF_X1 \o_values_reg[19][10]  (.D(o_values[10]), .CK(n_0_148), .Q(
      \o_values[19] [10]), .QN());
   DFF_X1 \o_values_reg[19][9]  (.D(o_values[9]), .CK(n_0_148), .Q(
      \o_values[19] [9]), .QN());
   DFF_X1 \o_values_reg[19][8]  (.D(o_values[8]), .CK(n_0_148), .Q(
      \o_values[19] [8]), .QN());
   DFF_X1 \o_values_reg[19][7]  (.D(o_values[7]), .CK(n_0_148), .Q(
      \o_values[19] [7]), .QN());
   DFF_X1 \o_values_reg[19][6]  (.D(o_values[6]), .CK(n_0_148), .Q(
      \o_values[19] [6]), .QN());
   DFF_X1 \o_values_reg[19][5]  (.D(o_values[5]), .CK(n_0_148), .Q(
      \o_values[19] [5]), .QN());
   DFF_X1 \o_values_reg[19][4]  (.D(o_values[4]), .CK(n_0_148), .Q(
      \o_values[19] [4]), .QN());
   DFF_X1 \o_values_reg[19][3]  (.D(o_values[3]), .CK(n_0_148), .Q(
      \o_values[19] [3]), .QN());
   DFF_X1 \o_values_reg[19][2]  (.D(o_values[2]), .CK(n_0_148), .Q(
      \o_values[19] [2]), .QN());
   DFF_X1 \o_values_reg[19][1]  (.D(o_values[1]), .CK(n_0_148), .Q(
      \o_values[19] [1]), .QN());
   DFF_X1 \o_values_reg[19][0]  (.D(o_values[0]), .CK(n_0_148), .Q(
      \o_values[19] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[18]_reg  (.CK(clk), .E(n_0_65), .SE(1'b0), 
      .GCK(n_0_149));
   DFF_X1 \o_values_reg[18][15]  (.D(o_values[15]), .CK(n_0_149), .Q(
      \o_values[18] [15]), .QN());
   DFF_X1 \o_values_reg[18][14]  (.D(o_values[14]), .CK(n_0_149), .Q(
      \o_values[18] [14]), .QN());
   DFF_X1 \o_values_reg[18][13]  (.D(o_values[13]), .CK(n_0_149), .Q(
      \o_values[18] [13]), .QN());
   DFF_X1 \o_values_reg[18][12]  (.D(o_values[12]), .CK(n_0_149), .Q(
      \o_values[18] [12]), .QN());
   DFF_X1 \o_values_reg[18][11]  (.D(o_values[11]), .CK(n_0_149), .Q(
      \o_values[18] [11]), .QN());
   DFF_X1 \o_values_reg[18][10]  (.D(o_values[10]), .CK(n_0_149), .Q(
      \o_values[18] [10]), .QN());
   DFF_X1 \o_values_reg[18][9]  (.D(o_values[9]), .CK(n_0_149), .Q(
      \o_values[18] [9]), .QN());
   DFF_X1 \o_values_reg[18][8]  (.D(o_values[8]), .CK(n_0_149), .Q(
      \o_values[18] [8]), .QN());
   DFF_X1 \o_values_reg[18][7]  (.D(o_values[7]), .CK(n_0_149), .Q(
      \o_values[18] [7]), .QN());
   DFF_X1 \o_values_reg[18][6]  (.D(o_values[6]), .CK(n_0_149), .Q(
      \o_values[18] [6]), .QN());
   DFF_X1 \o_values_reg[18][5]  (.D(o_values[5]), .CK(n_0_149), .Q(
      \o_values[18] [5]), .QN());
   DFF_X1 \o_values_reg[18][4]  (.D(o_values[4]), .CK(n_0_149), .Q(
      \o_values[18] [4]), .QN());
   DFF_X1 \o_values_reg[18][3]  (.D(o_values[3]), .CK(n_0_149), .Q(
      \o_values[18] [3]), .QN());
   DFF_X1 \o_values_reg[18][2]  (.D(o_values[2]), .CK(n_0_149), .Q(
      \o_values[18] [2]), .QN());
   DFF_X1 \o_values_reg[18][1]  (.D(o_values[1]), .CK(n_0_149), .Q(
      \o_values[18] [1]), .QN());
   DFF_X1 \o_values_reg[18][0]  (.D(o_values[0]), .CK(n_0_149), .Q(
      \o_values[18] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[17]_reg  (.CK(clk), .E(n_0_66), .SE(1'b0), 
      .GCK(n_0_150));
   DFF_X1 \o_values_reg[17][15]  (.D(o_values[15]), .CK(n_0_150), .Q(
      \o_values[17] [15]), .QN());
   DFF_X1 \o_values_reg[17][14]  (.D(o_values[14]), .CK(n_0_150), .Q(
      \o_values[17] [14]), .QN());
   DFF_X1 \o_values_reg[17][13]  (.D(o_values[13]), .CK(n_0_150), .Q(
      \o_values[17] [13]), .QN());
   DFF_X1 \o_values_reg[17][12]  (.D(o_values[12]), .CK(n_0_150), .Q(
      \o_values[17] [12]), .QN());
   DFF_X1 \o_values_reg[17][11]  (.D(o_values[11]), .CK(n_0_150), .Q(
      \o_values[17] [11]), .QN());
   DFF_X1 \o_values_reg[17][10]  (.D(o_values[10]), .CK(n_0_150), .Q(
      \o_values[17] [10]), .QN());
   DFF_X1 \o_values_reg[17][9]  (.D(o_values[9]), .CK(n_0_150), .Q(
      \o_values[17] [9]), .QN());
   DFF_X1 \o_values_reg[17][8]  (.D(o_values[8]), .CK(n_0_150), .Q(
      \o_values[17] [8]), .QN());
   DFF_X1 \o_values_reg[17][7]  (.D(o_values[7]), .CK(n_0_150), .Q(
      \o_values[17] [7]), .QN());
   DFF_X1 \o_values_reg[17][6]  (.D(o_values[6]), .CK(n_0_150), .Q(
      \o_values[17] [6]), .QN());
   DFF_X1 \o_values_reg[17][5]  (.D(o_values[5]), .CK(n_0_150), .Q(
      \o_values[17] [5]), .QN());
   DFF_X1 \o_values_reg[17][4]  (.D(o_values[4]), .CK(n_0_150), .Q(
      \o_values[17] [4]), .QN());
   DFF_X1 \o_values_reg[17][3]  (.D(o_values[3]), .CK(n_0_150), .Q(
      \o_values[17] [3]), .QN());
   DFF_X1 \o_values_reg[17][2]  (.D(o_values[2]), .CK(n_0_150), .Q(
      \o_values[17] [2]), .QN());
   DFF_X1 \o_values_reg[17][1]  (.D(o_values[1]), .CK(n_0_150), .Q(
      \o_values[17] [1]), .QN());
   DFF_X1 \o_values_reg[17][0]  (.D(o_values[0]), .CK(n_0_150), .Q(
      \o_values[17] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[16]_reg  (.CK(clk), .E(n_0_67), .SE(1'b0), 
      .GCK(n_0_151));
   DFF_X1 \o_values_reg[16][15]  (.D(o_values[15]), .CK(n_0_151), .Q(
      \o_values[16] [15]), .QN());
   DFF_X1 \o_values_reg[16][14]  (.D(o_values[14]), .CK(n_0_151), .Q(
      \o_values[16] [14]), .QN());
   DFF_X1 \o_values_reg[16][13]  (.D(o_values[13]), .CK(n_0_151), .Q(
      \o_values[16] [13]), .QN());
   DFF_X1 \o_values_reg[16][12]  (.D(o_values[12]), .CK(n_0_151), .Q(
      \o_values[16] [12]), .QN());
   DFF_X1 \o_values_reg[16][11]  (.D(o_values[11]), .CK(n_0_151), .Q(
      \o_values[16] [11]), .QN());
   DFF_X1 \o_values_reg[16][10]  (.D(o_values[10]), .CK(n_0_151), .Q(
      \o_values[16] [10]), .QN());
   DFF_X1 \o_values_reg[16][9]  (.D(o_values[9]), .CK(n_0_151), .Q(
      \o_values[16] [9]), .QN());
   DFF_X1 \o_values_reg[16][8]  (.D(o_values[8]), .CK(n_0_151), .Q(
      \o_values[16] [8]), .QN());
   DFF_X1 \o_values_reg[16][7]  (.D(o_values[7]), .CK(n_0_151), .Q(
      \o_values[16] [7]), .QN());
   DFF_X1 \o_values_reg[16][6]  (.D(o_values[6]), .CK(n_0_151), .Q(
      \o_values[16] [6]), .QN());
   DFF_X1 \o_values_reg[16][5]  (.D(o_values[5]), .CK(n_0_151), .Q(
      \o_values[16] [5]), .QN());
   DFF_X1 \o_values_reg[16][4]  (.D(o_values[4]), .CK(n_0_151), .Q(
      \o_values[16] [4]), .QN());
   DFF_X1 \o_values_reg[16][3]  (.D(o_values[3]), .CK(n_0_151), .Q(
      \o_values[16] [3]), .QN());
   DFF_X1 \o_values_reg[16][2]  (.D(o_values[2]), .CK(n_0_151), .Q(
      \o_values[16] [2]), .QN());
   DFF_X1 \o_values_reg[16][1]  (.D(o_values[1]), .CK(n_0_151), .Q(
      \o_values[16] [1]), .QN());
   DFF_X1 \o_values_reg[16][0]  (.D(o_values[0]), .CK(n_0_151), .Q(
      \o_values[16] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[15]_reg  (.CK(clk), .E(n_0_68), .SE(1'b0), 
      .GCK(n_0_152));
   DFF_X1 \o_values_reg[15][15]  (.D(o_values[15]), .CK(n_0_152), .Q(
      \o_values[15] [15]), .QN());
   DFF_X1 \o_values_reg[15][14]  (.D(o_values[14]), .CK(n_0_152), .Q(
      \o_values[15] [14]), .QN());
   DFF_X1 \o_values_reg[15][13]  (.D(o_values[13]), .CK(n_0_152), .Q(
      \o_values[15] [13]), .QN());
   DFF_X1 \o_values_reg[15][12]  (.D(o_values[12]), .CK(n_0_152), .Q(
      \o_values[15] [12]), .QN());
   DFF_X1 \o_values_reg[15][11]  (.D(o_values[11]), .CK(n_0_152), .Q(
      \o_values[15] [11]), .QN());
   DFF_X1 \o_values_reg[15][10]  (.D(o_values[10]), .CK(n_0_152), .Q(
      \o_values[15] [10]), .QN());
   DFF_X1 \o_values_reg[15][9]  (.D(o_values[9]), .CK(n_0_152), .Q(
      \o_values[15] [9]), .QN());
   DFF_X1 \o_values_reg[15][8]  (.D(o_values[8]), .CK(n_0_152), .Q(
      \o_values[15] [8]), .QN());
   DFF_X1 \o_values_reg[15][7]  (.D(o_values[7]), .CK(n_0_152), .Q(
      \o_values[15] [7]), .QN());
   DFF_X1 \o_values_reg[15][6]  (.D(o_values[6]), .CK(n_0_152), .Q(
      \o_values[15] [6]), .QN());
   DFF_X1 \o_values_reg[15][5]  (.D(o_values[5]), .CK(n_0_152), .Q(
      \o_values[15] [5]), .QN());
   DFF_X1 \o_values_reg[15][4]  (.D(o_values[4]), .CK(n_0_152), .Q(
      \o_values[15] [4]), .QN());
   DFF_X1 \o_values_reg[15][3]  (.D(o_values[3]), .CK(n_0_152), .Q(
      \o_values[15] [3]), .QN());
   DFF_X1 \o_values_reg[15][2]  (.D(o_values[2]), .CK(n_0_152), .Q(
      \o_values[15] [2]), .QN());
   DFF_X1 \o_values_reg[15][1]  (.D(o_values[1]), .CK(n_0_152), .Q(
      \o_values[15] [1]), .QN());
   DFF_X1 \o_values_reg[15][0]  (.D(o_values[0]), .CK(n_0_152), .Q(
      \o_values[15] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[14]_reg  (.CK(clk), .E(n_0_69), .SE(1'b0), 
      .GCK(n_0_153));
   DFF_X1 \o_values_reg[14][15]  (.D(o_values[15]), .CK(n_0_153), .Q(
      \o_values[14] [15]), .QN());
   DFF_X1 \o_values_reg[14][14]  (.D(o_values[14]), .CK(n_0_153), .Q(
      \o_values[14] [14]), .QN());
   DFF_X1 \o_values_reg[14][13]  (.D(o_values[13]), .CK(n_0_153), .Q(
      \o_values[14] [13]), .QN());
   DFF_X1 \o_values_reg[14][12]  (.D(o_values[12]), .CK(n_0_153), .Q(
      \o_values[14] [12]), .QN());
   DFF_X1 \o_values_reg[14][11]  (.D(o_values[11]), .CK(n_0_153), .Q(
      \o_values[14] [11]), .QN());
   DFF_X1 \o_values_reg[14][10]  (.D(o_values[10]), .CK(n_0_153), .Q(
      \o_values[14] [10]), .QN());
   DFF_X1 \o_values_reg[14][9]  (.D(o_values[9]), .CK(n_0_153), .Q(
      \o_values[14] [9]), .QN());
   DFF_X1 \o_values_reg[14][8]  (.D(o_values[8]), .CK(n_0_153), .Q(
      \o_values[14] [8]), .QN());
   DFF_X1 \o_values_reg[14][7]  (.D(o_values[7]), .CK(n_0_153), .Q(
      \o_values[14] [7]), .QN());
   DFF_X1 \o_values_reg[14][6]  (.D(o_values[6]), .CK(n_0_153), .Q(
      \o_values[14] [6]), .QN());
   DFF_X1 \o_values_reg[14][5]  (.D(o_values[5]), .CK(n_0_153), .Q(
      \o_values[14] [5]), .QN());
   DFF_X1 \o_values_reg[14][4]  (.D(o_values[4]), .CK(n_0_153), .Q(
      \o_values[14] [4]), .QN());
   DFF_X1 \o_values_reg[14][3]  (.D(o_values[3]), .CK(n_0_153), .Q(
      \o_values[14] [3]), .QN());
   DFF_X1 \o_values_reg[14][2]  (.D(o_values[2]), .CK(n_0_153), .Q(
      \o_values[14] [2]), .QN());
   DFF_X1 \o_values_reg[14][1]  (.D(o_values[1]), .CK(n_0_153), .Q(
      \o_values[14] [1]), .QN());
   DFF_X1 \o_values_reg[14][0]  (.D(o_values[0]), .CK(n_0_153), .Q(
      \o_values[14] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[13]_reg  (.CK(clk), .E(n_0_70), .SE(1'b0), 
      .GCK(n_0_154));
   DFF_X1 \o_values_reg[13][15]  (.D(o_values[15]), .CK(n_0_154), .Q(
      \o_values[13] [15]), .QN());
   DFF_X1 \o_values_reg[13][14]  (.D(o_values[14]), .CK(n_0_154), .Q(
      \o_values[13] [14]), .QN());
   DFF_X1 \o_values_reg[13][13]  (.D(o_values[13]), .CK(n_0_154), .Q(
      \o_values[13] [13]), .QN());
   DFF_X1 \o_values_reg[13][12]  (.D(o_values[12]), .CK(n_0_154), .Q(
      \o_values[13] [12]), .QN());
   DFF_X1 \o_values_reg[13][11]  (.D(o_values[11]), .CK(n_0_154), .Q(
      \o_values[13] [11]), .QN());
   DFF_X1 \o_values_reg[13][10]  (.D(o_values[10]), .CK(n_0_154), .Q(
      \o_values[13] [10]), .QN());
   DFF_X1 \o_values_reg[13][9]  (.D(o_values[9]), .CK(n_0_154), .Q(
      \o_values[13] [9]), .QN());
   DFF_X1 \o_values_reg[13][8]  (.D(o_values[8]), .CK(n_0_154), .Q(
      \o_values[13] [8]), .QN());
   DFF_X1 \o_values_reg[13][7]  (.D(o_values[7]), .CK(n_0_154), .Q(
      \o_values[13] [7]), .QN());
   DFF_X1 \o_values_reg[13][6]  (.D(o_values[6]), .CK(n_0_154), .Q(
      \o_values[13] [6]), .QN());
   DFF_X1 \o_values_reg[13][5]  (.D(o_values[5]), .CK(n_0_154), .Q(
      \o_values[13] [5]), .QN());
   DFF_X1 \o_values_reg[13][4]  (.D(o_values[4]), .CK(n_0_154), .Q(
      \o_values[13] [4]), .QN());
   DFF_X1 \o_values_reg[13][3]  (.D(o_values[3]), .CK(n_0_154), .Q(
      \o_values[13] [3]), .QN());
   DFF_X1 \o_values_reg[13][2]  (.D(o_values[2]), .CK(n_0_154), .Q(
      \o_values[13] [2]), .QN());
   DFF_X1 \o_values_reg[13][1]  (.D(o_values[1]), .CK(n_0_154), .Q(
      \o_values[13] [1]), .QN());
   DFF_X1 \o_values_reg[13][0]  (.D(o_values[0]), .CK(n_0_154), .Q(
      \o_values[13] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[12]_reg  (.CK(clk), .E(n_0_71), .SE(1'b0), 
      .GCK(n_0_155));
   DFF_X1 \o_values_reg[12][15]  (.D(o_values[15]), .CK(n_0_155), .Q(
      \o_values[12] [15]), .QN());
   DFF_X1 \o_values_reg[12][14]  (.D(o_values[14]), .CK(n_0_155), .Q(
      \o_values[12] [14]), .QN());
   DFF_X1 \o_values_reg[12][13]  (.D(o_values[13]), .CK(n_0_155), .Q(
      \o_values[12] [13]), .QN());
   DFF_X1 \o_values_reg[12][12]  (.D(o_values[12]), .CK(n_0_155), .Q(
      \o_values[12] [12]), .QN());
   DFF_X1 \o_values_reg[12][11]  (.D(o_values[11]), .CK(n_0_155), .Q(
      \o_values[12] [11]), .QN());
   DFF_X1 \o_values_reg[12][10]  (.D(o_values[10]), .CK(n_0_155), .Q(
      \o_values[12] [10]), .QN());
   DFF_X1 \o_values_reg[12][9]  (.D(o_values[9]), .CK(n_0_155), .Q(
      \o_values[12] [9]), .QN());
   DFF_X1 \o_values_reg[12][8]  (.D(o_values[8]), .CK(n_0_155), .Q(
      \o_values[12] [8]), .QN());
   DFF_X1 \o_values_reg[12][7]  (.D(o_values[7]), .CK(n_0_155), .Q(
      \o_values[12] [7]), .QN());
   DFF_X1 \o_values_reg[12][6]  (.D(o_values[6]), .CK(n_0_155), .Q(
      \o_values[12] [6]), .QN());
   DFF_X1 \o_values_reg[12][5]  (.D(o_values[5]), .CK(n_0_155), .Q(
      \o_values[12] [5]), .QN());
   DFF_X1 \o_values_reg[12][4]  (.D(o_values[4]), .CK(n_0_155), .Q(
      \o_values[12] [4]), .QN());
   DFF_X1 \o_values_reg[12][3]  (.D(o_values[3]), .CK(n_0_155), .Q(
      \o_values[12] [3]), .QN());
   DFF_X1 \o_values_reg[12][2]  (.D(o_values[2]), .CK(n_0_155), .Q(
      \o_values[12] [2]), .QN());
   DFF_X1 \o_values_reg[12][1]  (.D(o_values[1]), .CK(n_0_155), .Q(
      \o_values[12] [1]), .QN());
   DFF_X1 \o_values_reg[12][0]  (.D(o_values[0]), .CK(n_0_155), .Q(
      \o_values[12] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[11]_reg  (.CK(clk), .E(n_0_72), .SE(1'b0), 
      .GCK(n_0_156));
   DFF_X1 \o_values_reg[11][15]  (.D(o_values[15]), .CK(n_0_156), .Q(
      \o_values[11] [15]), .QN());
   DFF_X1 \o_values_reg[11][14]  (.D(o_values[14]), .CK(n_0_156), .Q(
      \o_values[11] [14]), .QN());
   DFF_X1 \o_values_reg[11][13]  (.D(o_values[13]), .CK(n_0_156), .Q(
      \o_values[11] [13]), .QN());
   DFF_X1 \o_values_reg[11][12]  (.D(o_values[12]), .CK(n_0_156), .Q(
      \o_values[11] [12]), .QN());
   DFF_X1 \o_values_reg[11][11]  (.D(o_values[11]), .CK(n_0_156), .Q(
      \o_values[11] [11]), .QN());
   DFF_X1 \o_values_reg[11][10]  (.D(o_values[10]), .CK(n_0_156), .Q(
      \o_values[11] [10]), .QN());
   DFF_X1 \o_values_reg[11][9]  (.D(o_values[9]), .CK(n_0_156), .Q(
      \o_values[11] [9]), .QN());
   DFF_X1 \o_values_reg[11][8]  (.D(o_values[8]), .CK(n_0_156), .Q(
      \o_values[11] [8]), .QN());
   DFF_X1 \o_values_reg[11][7]  (.D(o_values[7]), .CK(n_0_156), .Q(
      \o_values[11] [7]), .QN());
   DFF_X1 \o_values_reg[11][6]  (.D(o_values[6]), .CK(n_0_156), .Q(
      \o_values[11] [6]), .QN());
   DFF_X1 \o_values_reg[11][5]  (.D(o_values[5]), .CK(n_0_156), .Q(
      \o_values[11] [5]), .QN());
   DFF_X1 \o_values_reg[11][4]  (.D(o_values[4]), .CK(n_0_156), .Q(
      \o_values[11] [4]), .QN());
   DFF_X1 \o_values_reg[11][3]  (.D(o_values[3]), .CK(n_0_156), .Q(
      \o_values[11] [3]), .QN());
   DFF_X1 \o_values_reg[11][2]  (.D(o_values[2]), .CK(n_0_156), .Q(
      \o_values[11] [2]), .QN());
   DFF_X1 \o_values_reg[11][1]  (.D(o_values[1]), .CK(n_0_156), .Q(
      \o_values[11] [1]), .QN());
   DFF_X1 \o_values_reg[11][0]  (.D(o_values[0]), .CK(n_0_156), .Q(
      \o_values[11] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[10]_reg  (.CK(clk), .E(n_0_73), .SE(1'b0), 
      .GCK(n_0_157));
   DFF_X1 \o_values_reg[10][15]  (.D(o_values[15]), .CK(n_0_157), .Q(
      \o_values[10] [15]), .QN());
   DFF_X1 \o_values_reg[10][14]  (.D(o_values[14]), .CK(n_0_157), .Q(
      \o_values[10] [14]), .QN());
   DFF_X1 \o_values_reg[10][13]  (.D(o_values[13]), .CK(n_0_157), .Q(
      \o_values[10] [13]), .QN());
   DFF_X1 \o_values_reg[10][12]  (.D(o_values[12]), .CK(n_0_157), .Q(
      \o_values[10] [12]), .QN());
   DFF_X1 \o_values_reg[10][11]  (.D(o_values[11]), .CK(n_0_157), .Q(
      \o_values[10] [11]), .QN());
   DFF_X1 \o_values_reg[10][10]  (.D(o_values[10]), .CK(n_0_157), .Q(
      \o_values[10] [10]), .QN());
   DFF_X1 \o_values_reg[10][9]  (.D(o_values[9]), .CK(n_0_157), .Q(
      \o_values[10] [9]), .QN());
   DFF_X1 \o_values_reg[10][8]  (.D(o_values[8]), .CK(n_0_157), .Q(
      \o_values[10] [8]), .QN());
   DFF_X1 \o_values_reg[10][7]  (.D(o_values[7]), .CK(n_0_157), .Q(
      \o_values[10] [7]), .QN());
   DFF_X1 \o_values_reg[10][6]  (.D(o_values[6]), .CK(n_0_157), .Q(
      \o_values[10] [6]), .QN());
   DFF_X1 \o_values_reg[10][5]  (.D(o_values[5]), .CK(n_0_157), .Q(
      \o_values[10] [5]), .QN());
   DFF_X1 \o_values_reg[10][4]  (.D(o_values[4]), .CK(n_0_157), .Q(
      \o_values[10] [4]), .QN());
   DFF_X1 \o_values_reg[10][3]  (.D(o_values[3]), .CK(n_0_157), .Q(
      \o_values[10] [3]), .QN());
   DFF_X1 \o_values_reg[10][2]  (.D(o_values[2]), .CK(n_0_157), .Q(
      \o_values[10] [2]), .QN());
   DFF_X1 \o_values_reg[10][1]  (.D(o_values[1]), .CK(n_0_157), .Q(
      \o_values[10] [1]), .QN());
   DFF_X1 \o_values_reg[10][0]  (.D(o_values[0]), .CK(n_0_157), .Q(
      \o_values[10] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[9]_reg  (.CK(clk), .E(n_0_74), .SE(1'b0), 
      .GCK(n_0_158));
   DFF_X1 \o_values_reg[9][15]  (.D(o_values[15]), .CK(n_0_158), .Q(
      \o_values[9] [15]), .QN());
   DFF_X1 \o_values_reg[9][14]  (.D(o_values[14]), .CK(n_0_158), .Q(
      \o_values[9] [14]), .QN());
   DFF_X1 \o_values_reg[9][13]  (.D(o_values[13]), .CK(n_0_158), .Q(
      \o_values[9] [13]), .QN());
   DFF_X1 \o_values_reg[9][12]  (.D(o_values[12]), .CK(n_0_158), .Q(
      \o_values[9] [12]), .QN());
   DFF_X1 \o_values_reg[9][11]  (.D(o_values[11]), .CK(n_0_158), .Q(
      \o_values[9] [11]), .QN());
   DFF_X1 \o_values_reg[9][10]  (.D(o_values[10]), .CK(n_0_158), .Q(
      \o_values[9] [10]), .QN());
   DFF_X1 \o_values_reg[9][9]  (.D(o_values[9]), .CK(n_0_158), .Q(
      \o_values[9] [9]), .QN());
   DFF_X1 \o_values_reg[9][8]  (.D(o_values[8]), .CK(n_0_158), .Q(
      \o_values[9] [8]), .QN());
   DFF_X1 \o_values_reg[9][7]  (.D(o_values[7]), .CK(n_0_158), .Q(
      \o_values[9] [7]), .QN());
   DFF_X1 \o_values_reg[9][6]  (.D(o_values[6]), .CK(n_0_158), .Q(
      \o_values[9] [6]), .QN());
   DFF_X1 \o_values_reg[9][5]  (.D(o_values[5]), .CK(n_0_158), .Q(
      \o_values[9] [5]), .QN());
   DFF_X1 \o_values_reg[9][4]  (.D(o_values[4]), .CK(n_0_158), .Q(
      \o_values[9] [4]), .QN());
   DFF_X1 \o_values_reg[9][3]  (.D(o_values[3]), .CK(n_0_158), .Q(
      \o_values[9] [3]), .QN());
   DFF_X1 \o_values_reg[9][2]  (.D(o_values[2]), .CK(n_0_158), .Q(
      \o_values[9] [2]), .QN());
   DFF_X1 \o_values_reg[9][1]  (.D(o_values[1]), .CK(n_0_158), .Q(
      \o_values[9] [1]), .QN());
   DFF_X1 \o_values_reg[9][0]  (.D(o_values[0]), .CK(n_0_158), .Q(
      \o_values[9] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[8]_reg  (.CK(clk), .E(n_0_75), .SE(1'b0), 
      .GCK(n_0_159));
   DFF_X1 \o_values_reg[8][15]  (.D(o_values[15]), .CK(n_0_159), .Q(
      \o_values[8] [15]), .QN());
   DFF_X1 \o_values_reg[8][14]  (.D(o_values[14]), .CK(n_0_159), .Q(
      \o_values[8] [14]), .QN());
   DFF_X1 \o_values_reg[8][13]  (.D(o_values[13]), .CK(n_0_159), .Q(
      \o_values[8] [13]), .QN());
   DFF_X1 \o_values_reg[8][12]  (.D(o_values[12]), .CK(n_0_159), .Q(
      \o_values[8] [12]), .QN());
   DFF_X1 \o_values_reg[8][11]  (.D(o_values[11]), .CK(n_0_159), .Q(
      \o_values[8] [11]), .QN());
   DFF_X1 \o_values_reg[8][10]  (.D(o_values[10]), .CK(n_0_159), .Q(
      \o_values[8] [10]), .QN());
   DFF_X1 \o_values_reg[8][9]  (.D(o_values[9]), .CK(n_0_159), .Q(
      \o_values[8] [9]), .QN());
   DFF_X1 \o_values_reg[8][8]  (.D(o_values[8]), .CK(n_0_159), .Q(
      \o_values[8] [8]), .QN());
   DFF_X1 \o_values_reg[8][7]  (.D(o_values[7]), .CK(n_0_159), .Q(
      \o_values[8] [7]), .QN());
   DFF_X1 \o_values_reg[8][6]  (.D(o_values[6]), .CK(n_0_159), .Q(
      \o_values[8] [6]), .QN());
   DFF_X1 \o_values_reg[8][5]  (.D(o_values[5]), .CK(n_0_159), .Q(
      \o_values[8] [5]), .QN());
   DFF_X1 \o_values_reg[8][4]  (.D(o_values[4]), .CK(n_0_159), .Q(
      \o_values[8] [4]), .QN());
   DFF_X1 \o_values_reg[8][3]  (.D(o_values[3]), .CK(n_0_159), .Q(
      \o_values[8] [3]), .QN());
   DFF_X1 \o_values_reg[8][2]  (.D(o_values[2]), .CK(n_0_159), .Q(
      \o_values[8] [2]), .QN());
   DFF_X1 \o_values_reg[8][1]  (.D(o_values[1]), .CK(n_0_159), .Q(
      \o_values[8] [1]), .QN());
   DFF_X1 \o_values_reg[8][0]  (.D(o_values[0]), .CK(n_0_159), .Q(
      \o_values[8] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[7]_reg  (.CK(clk), .E(n_0_76), .SE(1'b0), 
      .GCK(n_0_160));
   DFF_X1 \o_values_reg[7][15]  (.D(o_values[15]), .CK(n_0_160), .Q(
      \o_values[7] [15]), .QN());
   DFF_X1 \o_values_reg[7][14]  (.D(o_values[14]), .CK(n_0_160), .Q(
      \o_values[7] [14]), .QN());
   DFF_X1 \o_values_reg[7][13]  (.D(o_values[13]), .CK(n_0_160), .Q(
      \o_values[7] [13]), .QN());
   DFF_X1 \o_values_reg[7][12]  (.D(o_values[12]), .CK(n_0_160), .Q(
      \o_values[7] [12]), .QN());
   DFF_X1 \o_values_reg[7][11]  (.D(o_values[11]), .CK(n_0_160), .Q(
      \o_values[7] [11]), .QN());
   DFF_X1 \o_values_reg[7][10]  (.D(o_values[10]), .CK(n_0_160), .Q(
      \o_values[7] [10]), .QN());
   DFF_X1 \o_values_reg[7][9]  (.D(o_values[9]), .CK(n_0_160), .Q(
      \o_values[7] [9]), .QN());
   DFF_X1 \o_values_reg[7][8]  (.D(o_values[8]), .CK(n_0_160), .Q(
      \o_values[7] [8]), .QN());
   DFF_X1 \o_values_reg[7][7]  (.D(o_values[7]), .CK(n_0_160), .Q(
      \o_values[7] [7]), .QN());
   DFF_X1 \o_values_reg[7][6]  (.D(o_values[6]), .CK(n_0_160), .Q(
      \o_values[7] [6]), .QN());
   DFF_X1 \o_values_reg[7][5]  (.D(o_values[5]), .CK(n_0_160), .Q(
      \o_values[7] [5]), .QN());
   DFF_X1 \o_values_reg[7][4]  (.D(o_values[4]), .CK(n_0_160), .Q(
      \o_values[7] [4]), .QN());
   DFF_X1 \o_values_reg[7][3]  (.D(o_values[3]), .CK(n_0_160), .Q(
      \o_values[7] [3]), .QN());
   DFF_X1 \o_values_reg[7][2]  (.D(o_values[2]), .CK(n_0_160), .Q(
      \o_values[7] [2]), .QN());
   DFF_X1 \o_values_reg[7][1]  (.D(o_values[1]), .CK(n_0_160), .Q(
      \o_values[7] [1]), .QN());
   DFF_X1 \o_values_reg[7][0]  (.D(o_values[0]), .CK(n_0_160), .Q(
      \o_values[7] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[6]_reg  (.CK(clk), .E(n_0_77), .SE(1'b0), 
      .GCK(n_0_161));
   DFF_X1 \o_values_reg[6][15]  (.D(o_values[15]), .CK(n_0_161), .Q(
      \o_values[6] [15]), .QN());
   DFF_X1 \o_values_reg[6][14]  (.D(o_values[14]), .CK(n_0_161), .Q(
      \o_values[6] [14]), .QN());
   DFF_X1 \o_values_reg[6][13]  (.D(o_values[13]), .CK(n_0_161), .Q(
      \o_values[6] [13]), .QN());
   DFF_X1 \o_values_reg[6][12]  (.D(o_values[12]), .CK(n_0_161), .Q(
      \o_values[6] [12]), .QN());
   DFF_X1 \o_values_reg[6][11]  (.D(o_values[11]), .CK(n_0_161), .Q(
      \o_values[6] [11]), .QN());
   DFF_X1 \o_values_reg[6][10]  (.D(o_values[10]), .CK(n_0_161), .Q(
      \o_values[6] [10]), .QN());
   DFF_X1 \o_values_reg[6][9]  (.D(o_values[9]), .CK(n_0_161), .Q(
      \o_values[6] [9]), .QN());
   DFF_X1 \o_values_reg[6][8]  (.D(o_values[8]), .CK(n_0_161), .Q(
      \o_values[6] [8]), .QN());
   DFF_X1 \o_values_reg[6][7]  (.D(o_values[7]), .CK(n_0_161), .Q(
      \o_values[6] [7]), .QN());
   DFF_X1 \o_values_reg[6][6]  (.D(o_values[6]), .CK(n_0_161), .Q(
      \o_values[6] [6]), .QN());
   DFF_X1 \o_values_reg[6][5]  (.D(o_values[5]), .CK(n_0_161), .Q(
      \o_values[6] [5]), .QN());
   DFF_X1 \o_values_reg[6][4]  (.D(o_values[4]), .CK(n_0_161), .Q(
      \o_values[6] [4]), .QN());
   DFF_X1 \o_values_reg[6][3]  (.D(o_values[3]), .CK(n_0_161), .Q(
      \o_values[6] [3]), .QN());
   DFF_X1 \o_values_reg[6][2]  (.D(o_values[2]), .CK(n_0_161), .Q(
      \o_values[6] [2]), .QN());
   DFF_X1 \o_values_reg[6][1]  (.D(o_values[1]), .CK(n_0_161), .Q(
      \o_values[6] [1]), .QN());
   DFF_X1 \o_values_reg[6][0]  (.D(o_values[0]), .CK(n_0_161), .Q(
      \o_values[6] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[5]_reg  (.CK(clk), .E(n_0_78), .SE(1'b0), 
      .GCK(n_0_162));
   DFF_X1 \o_values_reg[5][15]  (.D(o_values[15]), .CK(n_0_162), .Q(
      \o_values[5] [15]), .QN());
   DFF_X1 \o_values_reg[5][14]  (.D(o_values[14]), .CK(n_0_162), .Q(
      \o_values[5] [14]), .QN());
   DFF_X1 \o_values_reg[5][13]  (.D(o_values[13]), .CK(n_0_162), .Q(
      \o_values[5] [13]), .QN());
   DFF_X1 \o_values_reg[5][12]  (.D(o_values[12]), .CK(n_0_162), .Q(
      \o_values[5] [12]), .QN());
   DFF_X1 \o_values_reg[5][11]  (.D(o_values[11]), .CK(n_0_162), .Q(
      \o_values[5] [11]), .QN());
   DFF_X1 \o_values_reg[5][10]  (.D(o_values[10]), .CK(n_0_162), .Q(
      \o_values[5] [10]), .QN());
   DFF_X1 \o_values_reg[5][9]  (.D(o_values[9]), .CK(n_0_162), .Q(
      \o_values[5] [9]), .QN());
   DFF_X1 \o_values_reg[5][8]  (.D(o_values[8]), .CK(n_0_162), .Q(
      \o_values[5] [8]), .QN());
   DFF_X1 \o_values_reg[5][7]  (.D(o_values[7]), .CK(n_0_162), .Q(
      \o_values[5] [7]), .QN());
   DFF_X1 \o_values_reg[5][6]  (.D(o_values[6]), .CK(n_0_162), .Q(
      \o_values[5] [6]), .QN());
   DFF_X1 \o_values_reg[5][5]  (.D(o_values[5]), .CK(n_0_162), .Q(
      \o_values[5] [5]), .QN());
   DFF_X1 \o_values_reg[5][4]  (.D(o_values[4]), .CK(n_0_162), .Q(
      \o_values[5] [4]), .QN());
   DFF_X1 \o_values_reg[5][3]  (.D(o_values[3]), .CK(n_0_162), .Q(
      \o_values[5] [3]), .QN());
   DFF_X1 \o_values_reg[5][2]  (.D(o_values[2]), .CK(n_0_162), .Q(
      \o_values[5] [2]), .QN());
   DFF_X1 \o_values_reg[5][1]  (.D(o_values[1]), .CK(n_0_162), .Q(
      \o_values[5] [1]), .QN());
   DFF_X1 \o_values_reg[5][0]  (.D(o_values[0]), .CK(n_0_162), .Q(
      \o_values[5] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[4]_reg  (.CK(clk), .E(n_0_79), .SE(1'b0), 
      .GCK(n_0_163));
   DFF_X1 \o_values_reg[4][15]  (.D(o_values[15]), .CK(n_0_163), .Q(
      \o_values[4] [15]), .QN());
   DFF_X1 \o_values_reg[4][14]  (.D(o_values[14]), .CK(n_0_163), .Q(
      \o_values[4] [14]), .QN());
   DFF_X1 \o_values_reg[4][13]  (.D(o_values[13]), .CK(n_0_163), .Q(
      \o_values[4] [13]), .QN());
   DFF_X1 \o_values_reg[4][12]  (.D(o_values[12]), .CK(n_0_163), .Q(
      \o_values[4] [12]), .QN());
   DFF_X1 \o_values_reg[4][11]  (.D(o_values[11]), .CK(n_0_163), .Q(
      \o_values[4] [11]), .QN());
   DFF_X1 \o_values_reg[4][10]  (.D(o_values[10]), .CK(n_0_163), .Q(
      \o_values[4] [10]), .QN());
   DFF_X1 \o_values_reg[4][9]  (.D(o_values[9]), .CK(n_0_163), .Q(
      \o_values[4] [9]), .QN());
   DFF_X1 \o_values_reg[4][8]  (.D(o_values[8]), .CK(n_0_163), .Q(
      \o_values[4] [8]), .QN());
   DFF_X1 \o_values_reg[4][7]  (.D(o_values[7]), .CK(n_0_163), .Q(
      \o_values[4] [7]), .QN());
   DFF_X1 \o_values_reg[4][6]  (.D(o_values[6]), .CK(n_0_163), .Q(
      \o_values[4] [6]), .QN());
   DFF_X1 \o_values_reg[4][5]  (.D(o_values[5]), .CK(n_0_163), .Q(
      \o_values[4] [5]), .QN());
   DFF_X1 \o_values_reg[4][4]  (.D(o_values[4]), .CK(n_0_163), .Q(
      \o_values[4] [4]), .QN());
   DFF_X1 \o_values_reg[4][3]  (.D(o_values[3]), .CK(n_0_163), .Q(
      \o_values[4] [3]), .QN());
   DFF_X1 \o_values_reg[4][2]  (.D(o_values[2]), .CK(n_0_163), .Q(
      \o_values[4] [2]), .QN());
   DFF_X1 \o_values_reg[4][1]  (.D(o_values[1]), .CK(n_0_163), .Q(
      \o_values[4] [1]), .QN());
   DFF_X1 \o_values_reg[4][0]  (.D(o_values[0]), .CK(n_0_163), .Q(
      \o_values[4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[3]_reg  (.CK(clk), .E(n_0_80), .SE(1'b0), 
      .GCK(n_0_164));
   DFF_X1 \o_values_reg[3][15]  (.D(o_values[15]), .CK(n_0_164), .Q(
      \o_values[3] [15]), .QN());
   DFF_X1 \o_values_reg[3][14]  (.D(o_values[14]), .CK(n_0_164), .Q(
      \o_values[3] [14]), .QN());
   DFF_X1 \o_values_reg[3][13]  (.D(o_values[13]), .CK(n_0_164), .Q(
      \o_values[3] [13]), .QN());
   DFF_X1 \o_values_reg[3][12]  (.D(o_values[12]), .CK(n_0_164), .Q(
      \o_values[3] [12]), .QN());
   DFF_X1 \o_values_reg[3][11]  (.D(o_values[11]), .CK(n_0_164), .Q(
      \o_values[3] [11]), .QN());
   DFF_X1 \o_values_reg[3][10]  (.D(o_values[10]), .CK(n_0_164), .Q(
      \o_values[3] [10]), .QN());
   DFF_X1 \o_values_reg[3][9]  (.D(o_values[9]), .CK(n_0_164), .Q(
      \o_values[3] [9]), .QN());
   DFF_X1 \o_values_reg[3][8]  (.D(o_values[8]), .CK(n_0_164), .Q(
      \o_values[3] [8]), .QN());
   DFF_X1 \o_values_reg[3][7]  (.D(o_values[7]), .CK(n_0_164), .Q(
      \o_values[3] [7]), .QN());
   DFF_X1 \o_values_reg[3][6]  (.D(o_values[6]), .CK(n_0_164), .Q(
      \o_values[3] [6]), .QN());
   DFF_X1 \o_values_reg[3][5]  (.D(o_values[5]), .CK(n_0_164), .Q(
      \o_values[3] [5]), .QN());
   DFF_X1 \o_values_reg[3][4]  (.D(o_values[4]), .CK(n_0_164), .Q(
      \o_values[3] [4]), .QN());
   DFF_X1 \o_values_reg[3][3]  (.D(o_values[3]), .CK(n_0_164), .Q(
      \o_values[3] [3]), .QN());
   DFF_X1 \o_values_reg[3][2]  (.D(o_values[2]), .CK(n_0_164), .Q(
      \o_values[3] [2]), .QN());
   DFF_X1 \o_values_reg[3][1]  (.D(o_values[1]), .CK(n_0_164), .Q(
      \o_values[3] [1]), .QN());
   DFF_X1 \o_values_reg[3][0]  (.D(o_values[0]), .CK(n_0_164), .Q(
      \o_values[3] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[2]_reg  (.CK(clk), .E(n_0_81), .SE(1'b0), 
      .GCK(n_0_165));
   DFF_X1 \o_values_reg[2][15]  (.D(o_values[15]), .CK(n_0_165), .Q(
      \o_values[2] [15]), .QN());
   DFF_X1 \o_values_reg[2][14]  (.D(o_values[14]), .CK(n_0_165), .Q(
      \o_values[2] [14]), .QN());
   DFF_X1 \o_values_reg[2][13]  (.D(o_values[13]), .CK(n_0_165), .Q(
      \o_values[2] [13]), .QN());
   DFF_X1 \o_values_reg[2][12]  (.D(o_values[12]), .CK(n_0_165), .Q(
      \o_values[2] [12]), .QN());
   DFF_X1 \o_values_reg[2][11]  (.D(o_values[11]), .CK(n_0_165), .Q(
      \o_values[2] [11]), .QN());
   DFF_X1 \o_values_reg[2][10]  (.D(o_values[10]), .CK(n_0_165), .Q(
      \o_values[2] [10]), .QN());
   DFF_X1 \o_values_reg[2][9]  (.D(o_values[9]), .CK(n_0_165), .Q(
      \o_values[2] [9]), .QN());
   DFF_X1 \o_values_reg[2][8]  (.D(o_values[8]), .CK(n_0_165), .Q(
      \o_values[2] [8]), .QN());
   DFF_X1 \o_values_reg[2][7]  (.D(o_values[7]), .CK(n_0_165), .Q(
      \o_values[2] [7]), .QN());
   DFF_X1 \o_values_reg[2][6]  (.D(o_values[6]), .CK(n_0_165), .Q(
      \o_values[2] [6]), .QN());
   DFF_X1 \o_values_reg[2][5]  (.D(o_values[5]), .CK(n_0_165), .Q(
      \o_values[2] [5]), .QN());
   DFF_X1 \o_values_reg[2][4]  (.D(o_values[4]), .CK(n_0_165), .Q(
      \o_values[2] [4]), .QN());
   DFF_X1 \o_values_reg[2][3]  (.D(o_values[3]), .CK(n_0_165), .Q(
      \o_values[2] [3]), .QN());
   DFF_X1 \o_values_reg[2][2]  (.D(o_values[2]), .CK(n_0_165), .Q(
      \o_values[2] [2]), .QN());
   DFF_X1 \o_values_reg[2][1]  (.D(o_values[1]), .CK(n_0_165), .Q(
      \o_values[2] [1]), .QN());
   DFF_X1 \o_values_reg[2][0]  (.D(o_values[0]), .CK(n_0_165), .Q(
      \o_values[2] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[1]_reg  (.CK(clk), .E(n_0_82), .SE(1'b0), 
      .GCK(n_0_166));
   DFF_X1 \o_values_reg[1][15]  (.D(o_values[15]), .CK(n_0_166), .Q(
      \o_values[1] [15]), .QN());
   DFF_X1 \o_values_reg[1][14]  (.D(o_values[14]), .CK(n_0_166), .Q(
      \o_values[1] [14]), .QN());
   DFF_X1 \o_values_reg[1][13]  (.D(o_values[13]), .CK(n_0_166), .Q(
      \o_values[1] [13]), .QN());
   DFF_X1 \o_values_reg[1][12]  (.D(o_values[12]), .CK(n_0_166), .Q(
      \o_values[1] [12]), .QN());
   DFF_X1 \o_values_reg[1][11]  (.D(o_values[11]), .CK(n_0_166), .Q(
      \o_values[1] [11]), .QN());
   DFF_X1 \o_values_reg[1][10]  (.D(o_values[10]), .CK(n_0_166), .Q(
      \o_values[1] [10]), .QN());
   DFF_X1 \o_values_reg[1][9]  (.D(o_values[9]), .CK(n_0_166), .Q(
      \o_values[1] [9]), .QN());
   DFF_X1 \o_values_reg[1][8]  (.D(o_values[8]), .CK(n_0_166), .Q(
      \o_values[1] [8]), .QN());
   DFF_X1 \o_values_reg[1][7]  (.D(o_values[7]), .CK(n_0_166), .Q(
      \o_values[1] [7]), .QN());
   DFF_X1 \o_values_reg[1][6]  (.D(o_values[6]), .CK(n_0_166), .Q(
      \o_values[1] [6]), .QN());
   DFF_X1 \o_values_reg[1][5]  (.D(o_values[5]), .CK(n_0_166), .Q(
      \o_values[1] [5]), .QN());
   DFF_X1 \o_values_reg[1][4]  (.D(o_values[4]), .CK(n_0_166), .Q(
      \o_values[1] [4]), .QN());
   DFF_X1 \o_values_reg[1][3]  (.D(o_values[3]), .CK(n_0_166), .Q(
      \o_values[1] [3]), .QN());
   DFF_X1 \o_values_reg[1][2]  (.D(o_values[2]), .CK(n_0_166), .Q(
      \o_values[1] [2]), .QN());
   DFF_X1 \o_values_reg[1][1]  (.D(o_values[1]), .CK(n_0_166), .Q(
      \o_values[1] [1]), .QN());
   DFF_X1 \o_values_reg[1][0]  (.D(o_values[0]), .CK(n_0_166), .Q(
      \o_values[1] [0]), .QN());
   CLKGATETST_X1 \clk_gate_o_values_reg[0]_reg  (.CK(clk), .E(n_0_83), .SE(1'b0), 
      .GCK(n_0_167));
   DFF_X1 \o_values_reg[0][15]  (.D(o_values[15]), .CK(n_0_167), .Q(
      \o_values[0] [15]), .QN());
   DFF_X1 \o_values_reg[0][14]  (.D(o_values[14]), .CK(n_0_167), .Q(
      \o_values[0] [14]), .QN());
   DFF_X1 \o_values_reg[0][13]  (.D(o_values[13]), .CK(n_0_167), .Q(
      \o_values[0] [13]), .QN());
   DFF_X1 \o_values_reg[0][12]  (.D(o_values[12]), .CK(n_0_167), .Q(
      \o_values[0] [12]), .QN());
   DFF_X1 \o_values_reg[0][11]  (.D(o_values[11]), .CK(n_0_167), .Q(
      \o_values[0] [11]), .QN());
   DFF_X1 \o_values_reg[0][10]  (.D(o_values[10]), .CK(n_0_167), .Q(
      \o_values[0] [10]), .QN());
   DFF_X1 \o_values_reg[0][9]  (.D(o_values[9]), .CK(n_0_167), .Q(
      \o_values[0] [9]), .QN());
   DFF_X1 \o_values_reg[0][8]  (.D(o_values[8]), .CK(n_0_167), .Q(
      \o_values[0] [8]), .QN());
   DFF_X1 \o_values_reg[0][7]  (.D(o_values[7]), .CK(n_0_167), .Q(
      \o_values[0] [7]), .QN());
   DFF_X1 \o_values_reg[0][6]  (.D(o_values[6]), .CK(n_0_167), .Q(
      \o_values[0] [6]), .QN());
   DFF_X1 \o_values_reg[0][5]  (.D(o_values[5]), .CK(n_0_167), .Q(
      \o_values[0] [5]), .QN());
   DFF_X1 \o_values_reg[0][4]  (.D(o_values[4]), .CK(n_0_167), .Q(
      \o_values[0] [4]), .QN());
   DFF_X1 \o_values_reg[0][3]  (.D(o_values[3]), .CK(n_0_167), .Q(
      \o_values[0] [3]), .QN());
   DFF_X1 \o_values_reg[0][2]  (.D(o_values[2]), .CK(n_0_167), .Q(
      \o_values[0] [2]), .QN());
   DFF_X1 \o_values_reg[0][1]  (.D(o_values[1]), .CK(n_0_167), .Q(
      \o_values[0] [1]), .QN());
   DFF_X1 \o_values_reg[0][0]  (.D(o_values[0]), .CK(n_0_167), .Q(
      \o_values[0] [0]), .QN());
   AND2_X1 i_0_0_0 (.A1(n_0_0_52), .A2(load_value[0]), .ZN(o_values[0]));
   AND2_X1 i_0_0_1 (.A1(n_0_0_52), .A2(load_value[1]), .ZN(o_values[1]));
   AND2_X1 i_0_0_2 (.A1(n_0_0_52), .A2(load_value[2]), .ZN(o_values[2]));
   AND2_X1 i_0_0_3 (.A1(n_0_0_52), .A2(load_value[3]), .ZN(o_values[3]));
   AND2_X1 i_0_0_4 (.A1(n_0_0_52), .A2(load_value[4]), .ZN(o_values[4]));
   AND2_X1 i_0_0_5 (.A1(n_0_0_52), .A2(load_value[5]), .ZN(o_values[5]));
   AND2_X1 i_0_0_6 (.A1(n_0_0_52), .A2(load_value[6]), .ZN(o_values[6]));
   AND2_X1 i_0_0_7 (.A1(n_0_0_52), .A2(load_value[7]), .ZN(o_values[7]));
   AND2_X1 i_0_0_8 (.A1(n_0_0_52), .A2(load_value[8]), .ZN(o_values[8]));
   AND2_X1 i_0_0_9 (.A1(n_0_0_52), .A2(load_value[9]), .ZN(o_values[9]));
   AND2_X1 i_0_0_10 (.A1(n_0_0_52), .A2(load_value[10]), .ZN(o_values[10]));
   AND2_X1 i_0_0_11 (.A1(n_0_0_52), .A2(load_value[11]), .ZN(o_values[11]));
   AND2_X1 i_0_0_12 (.A1(n_0_0_52), .A2(load_value[12]), .ZN(o_values[12]));
   AND2_X1 i_0_0_13 (.A1(n_0_0_52), .A2(load_value[13]), .ZN(o_values[13]));
   AND2_X1 i_0_0_14 (.A1(n_0_0_52), .A2(load_value[14]), .ZN(o_values[14]));
   AND2_X1 i_0_0_15 (.A1(n_0_0_52), .A2(load_value[15]), .ZN(o_values[15]));
   OAI21_X1 i_0_0_16 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_0), .ZN(n_0_83));
   OAI21_X1 i_0_0_17 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_0), .ZN(n_0_82));
   OAI21_X1 i_0_0_18 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_0), .ZN(n_0_81));
   OAI21_X1 i_0_0_19 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_0), .ZN(n_0_80));
   NAND2_X1 i_0_0_20 (.A1(n_0_0_42), .A2(n_0_0_30), .ZN(n_0_0_0));
   OAI21_X1 i_0_0_21 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_1), .ZN(n_0_79));
   OAI21_X1 i_0_0_22 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_1), .ZN(n_0_78));
   OAI21_X1 i_0_0_23 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_1), .ZN(n_0_77));
   OAI21_X1 i_0_0_24 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_1), .ZN(n_0_76));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_30), .A2(n_0_0_22), .ZN(n_0_0_1));
   OAI21_X1 i_0_0_26 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_2), .ZN(n_0_75));
   OAI21_X1 i_0_0_27 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_2), .ZN(n_0_74));
   OAI21_X1 i_0_0_28 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_2), .ZN(n_0_73));
   OAI21_X1 i_0_0_29 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_2), .ZN(n_0_72));
   NAND2_X1 i_0_0_30 (.A1(n_0_0_30), .A2(n_0_0_24), .ZN(n_0_0_2));
   OAI21_X1 i_0_0_31 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_3), .ZN(n_0_71));
   OAI21_X1 i_0_0_32 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_3), .ZN(n_0_70));
   OAI21_X1 i_0_0_33 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_3), .ZN(n_0_69));
   OAI21_X1 i_0_0_34 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_3), .ZN(n_0_68));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_32), .A2(n_0_0_30), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_36 (.A(n_0_0_52), .B1(n_0_0_39), .B2(n_0_0_15), .ZN(n_0_67));
   OAI21_X1 i_0_0_37 (.A(n_0_0_52), .B1(n_0_0_39), .B2(n_0_0_16), .ZN(n_0_66));
   OAI21_X1 i_0_0_38 (.A(n_0_0_52), .B1(n_0_0_39), .B2(n_0_0_17), .ZN(n_0_65));
   OAI21_X1 i_0_0_39 (.A(n_0_0_52), .B1(n_0_0_39), .B2(n_0_0_18), .ZN(n_0_64));
   OAI21_X1 i_0_0_40 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_4), .ZN(n_0_63));
   OAI21_X1 i_0_0_41 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_4), .ZN(n_0_62));
   OAI21_X1 i_0_0_42 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_4), .ZN(n_0_61));
   OAI21_X1 i_0_0_43 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_4), .ZN(n_0_60));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_40), .A2(n_0_0_22), .ZN(n_0_0_4));
   OAI21_X1 i_0_0_45 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_5), .ZN(n_0_59));
   OAI21_X1 i_0_0_46 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_5), .ZN(n_0_58));
   OAI21_X1 i_0_0_47 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_5), .ZN(n_0_57));
   OAI21_X1 i_0_0_48 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_5), .ZN(n_0_56));
   NAND2_X1 i_0_0_49 (.A1(n_0_0_40), .A2(n_0_0_24), .ZN(n_0_0_5));
   OAI21_X1 i_0_0_50 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_6), .ZN(n_0_55));
   OAI21_X1 i_0_0_51 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_6), .ZN(n_0_54));
   OAI21_X1 i_0_0_52 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_6), .ZN(n_0_53));
   OAI21_X1 i_0_0_53 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_6), .ZN(n_0_52));
   NAND2_X1 i_0_0_54 (.A1(n_0_0_40), .A2(n_0_0_32), .ZN(n_0_0_6));
   OAI21_X1 i_0_0_55 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_7), .ZN(n_0_51));
   OAI21_X1 i_0_0_56 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_7), .ZN(n_0_50));
   OAI21_X1 i_0_0_57 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_7), .ZN(n_0_49));
   OAI21_X1 i_0_0_58 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_7), .ZN(n_0_48));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_42), .A2(n_0_0_11), .ZN(n_0_0_7));
   OAI21_X1 i_0_0_60 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_8), .ZN(n_0_47));
   OAI21_X1 i_0_0_61 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_8), .ZN(n_0_46));
   OAI21_X1 i_0_0_62 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_8), .ZN(n_0_45));
   OAI21_X1 i_0_0_63 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_8), .ZN(n_0_44));
   NAND2_X1 i_0_0_64 (.A1(n_0_0_22), .A2(n_0_0_11), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_65 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_9), .ZN(n_0_43));
   OAI21_X1 i_0_0_66 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_9), .ZN(n_0_42));
   OAI21_X1 i_0_0_67 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_9), .ZN(n_0_41));
   OAI21_X1 i_0_0_68 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_9), .ZN(n_0_40));
   NAND2_X1 i_0_0_69 (.A1(n_0_0_24), .A2(n_0_0_11), .ZN(n_0_0_9));
   OAI21_X1 i_0_0_70 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_10), .ZN(n_0_39));
   OAI21_X1 i_0_0_71 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_10), .ZN(n_0_38));
   OAI21_X1 i_0_0_72 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_10), .ZN(n_0_37));
   OAI21_X1 i_0_0_73 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_10), .ZN(n_0_36));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_32), .A2(n_0_0_11), .ZN(n_0_0_10));
   AND2_X1 i_0_0_75 (.A1(n_0_0_50), .A2(load_address[5]), .ZN(n_0_0_11));
   OAI21_X1 i_0_0_76 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_12), .ZN(n_0_35));
   OAI21_X1 i_0_0_77 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_12), .ZN(n_0_34));
   OAI21_X1 i_0_0_78 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_12), .ZN(n_0_33));
   OAI21_X1 i_0_0_79 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_12), .ZN(n_0_32));
   NAND3_X1 i_0_0_80 (.A1(load_address[5]), .A2(load_address[4]), .A3(n_0_0_42), 
      .ZN(n_0_0_12));
   OAI21_X1 i_0_0_81 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_13), .ZN(n_0_31));
   OAI21_X1 i_0_0_82 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_13), .ZN(n_0_30));
   OAI21_X1 i_0_0_83 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_13), .ZN(n_0_29));
   OAI21_X1 i_0_0_84 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_13), .ZN(n_0_28));
   NAND3_X1 i_0_0_85 (.A1(load_address[5]), .A2(load_address[4]), .A3(n_0_0_22), 
      .ZN(n_0_0_13));
   OAI21_X1 i_0_0_86 (.A(n_0_0_52), .B1(n_0_0_15), .B2(n_0_0_14), .ZN(n_0_27));
   OAI21_X1 i_0_0_87 (.A(n_0_0_52), .B1(n_0_0_16), .B2(n_0_0_14), .ZN(n_0_26));
   OAI21_X1 i_0_0_88 (.A(n_0_0_52), .B1(n_0_0_17), .B2(n_0_0_14), .ZN(n_0_25));
   OAI21_X1 i_0_0_89 (.A(n_0_0_52), .B1(n_0_0_18), .B2(n_0_0_14), .ZN(n_0_24));
   NAND3_X1 i_0_0_90 (.A1(load_address[5]), .A2(load_address[4]), .A3(n_0_0_24), 
      .ZN(n_0_0_14));
   OAI21_X1 i_0_0_91 (.A(n_0_0_52), .B1(n_0_0_20), .B2(n_0_0_15), .ZN(n_0_23));
   NAND3_X1 i_0_0_92 (.A1(n_0_0_19), .A2(n_0_0_46), .A3(n_0_0_47), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_93 (.A(n_0_0_52), .B1(n_0_0_20), .B2(n_0_0_16), .ZN(n_0_22));
   NAND3_X1 i_0_0_94 (.A1(n_0_0_19), .A2(n_0_0_47), .A3(load_address[0]), 
      .ZN(n_0_0_16));
   OAI21_X1 i_0_0_95 (.A(n_0_0_52), .B1(n_0_0_20), .B2(n_0_0_17), .ZN(n_0_21));
   NAND3_X1 i_0_0_96 (.A1(load_address[1]), .A2(n_0_0_19), .A3(n_0_0_46), 
      .ZN(n_0_0_17));
   OAI21_X1 i_0_0_97 (.A(n_0_0_52), .B1(n_0_0_20), .B2(n_0_0_18), .ZN(n_0_20));
   NAND3_X1 i_0_0_98 (.A1(load_address[1]), .A2(load_address[0]), .A3(n_0_0_19), 
      .ZN(n_0_0_18));
   NOR2_X1 i_0_0_99 (.A1(n_0_0_37), .A2(load_address[6]), .ZN(n_0_0_19));
   NAND3_X1 i_0_0_100 (.A1(load_address[5]), .A2(load_address[4]), .A3(n_0_0_32), 
      .ZN(n_0_0_20));
   OAI21_X1 i_0_0_101 (.A(n_0_0_52), .B1(n_0_0_41), .B2(n_0_0_25), .ZN(n_0_19));
   OAI21_X1 i_0_0_102 (.A(n_0_0_52), .B1(n_0_0_41), .B2(n_0_0_26), .ZN(n_0_18));
   OAI21_X1 i_0_0_103 (.A(n_0_0_52), .B1(n_0_0_41), .B2(n_0_0_27), .ZN(n_0_17));
   OAI21_X1 i_0_0_104 (.A(n_0_0_52), .B1(n_0_0_41), .B2(n_0_0_28), .ZN(n_0_16));
   OAI21_X1 i_0_0_105 (.A(n_0_0_52), .B1(n_0_0_25), .B2(n_0_0_21), .ZN(n_0_15));
   OAI21_X1 i_0_0_106 (.A(n_0_0_52), .B1(n_0_0_26), .B2(n_0_0_21), .ZN(n_0_14));
   OAI21_X1 i_0_0_107 (.A(n_0_0_52), .B1(n_0_0_27), .B2(n_0_0_21), .ZN(n_0_13));
   OAI21_X1 i_0_0_108 (.A(n_0_0_52), .B1(n_0_0_28), .B2(n_0_0_21), .ZN(n_0_12));
   NAND2_X1 i_0_0_109 (.A1(n_0_0_49), .A2(load_address[2]), .ZN(n_0_0_21));
   NOR2_X1 i_0_0_110 (.A1(n_0_0_48), .A2(load_address[3]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_111 (.A(n_0_0_52), .B1(n_0_0_25), .B2(n_0_0_23), .ZN(n_0_11));
   OAI21_X1 i_0_0_112 (.A(n_0_0_52), .B1(n_0_0_26), .B2(n_0_0_23), .ZN(n_0_10));
   OAI21_X1 i_0_0_113 (.A(n_0_0_52), .B1(n_0_0_27), .B2(n_0_0_23), .ZN(n_0_9));
   OAI21_X1 i_0_0_114 (.A(n_0_0_52), .B1(n_0_0_28), .B2(n_0_0_23), .ZN(n_0_8));
   NAND2_X1 i_0_0_115 (.A1(n_0_0_48), .A2(load_address[3]), .ZN(n_0_0_23));
   NOR2_X1 i_0_0_116 (.A1(n_0_0_49), .A2(load_address[2]), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_117 (.A(n_0_0_52), .B1(n_0_0_31), .B2(n_0_0_25), .ZN(n_0_7));
   OR2_X1 i_0_0_118 (.A1(n_0_0_33), .A2(n_0_0_29), .ZN(n_0_0_25));
   OAI21_X1 i_0_0_119 (.A(n_0_0_52), .B1(n_0_0_31), .B2(n_0_0_26), .ZN(n_0_6));
   OR2_X1 i_0_0_120 (.A1(n_0_0_34), .A2(n_0_0_29), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_121 (.A(n_0_0_52), .B1(n_0_0_31), .B2(n_0_0_27), .ZN(n_0_5));
   OR2_X1 i_0_0_122 (.A1(n_0_0_35), .A2(n_0_0_29), .ZN(n_0_0_27));
   OAI21_X1 i_0_0_123 (.A(n_0_0_52), .B1(n_0_0_31), .B2(n_0_0_28), .ZN(n_0_4));
   OR2_X1 i_0_0_124 (.A1(n_0_0_45), .A2(n_0_0_29), .ZN(n_0_0_28));
   NAND3_X1 i_0_0_125 (.A1(load_address[6]), .A2(n_0_0_38), .A3(n_0_0_30), 
      .ZN(n_0_0_29));
   NOR2_X1 i_0_0_126 (.A1(load_address[5]), .A2(load_address[4]), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_127 (.A1(load_address[3]), .A2(load_address[2]), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_128 (.A1(n_0_0_49), .A2(n_0_0_48), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_129 (.A(n_0_0_52), .B1(n_0_0_36), .B2(n_0_0_33), .ZN(n_0_3));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_47), .A2(n_0_0_46), .ZN(n_0_0_33));
   OAI21_X1 i_0_0_131 (.A(n_0_0_52), .B1(n_0_0_36), .B2(n_0_0_34), .ZN(n_0_2));
   NAND2_X1 i_0_0_132 (.A1(n_0_0_47), .A2(load_address[0]), .ZN(n_0_0_34));
   OAI21_X1 i_0_0_133 (.A(n_0_0_52), .B1(n_0_0_36), .B2(n_0_0_35), .ZN(n_0_1));
   NAND2_X1 i_0_0_134 (.A1(n_0_0_46), .A2(load_address[1]), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_135 (.A(n_0_0_52), .B1(n_0_0_45), .B2(n_0_0_36), .ZN(n_0_0));
   NAND4_X1 i_0_0_136 (.A1(load_address[6]), .A2(n_0_0_42), .A3(n_0_0_40), 
      .A4(n_0_0_38), .ZN(n_0_0_36));
   INV_X1 i_0_0_137 (.A(n_0_0_38), .ZN(n_0_0_37));
   NOR4_X1 i_0_0_138 (.A1(n_0_0_44), .A2(n_0_0_43), .A3(load_address[8]), 
      .A4(load_address[7]), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_42), .A2(n_0_0_40), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_140 (.A1(n_0_0_50), .A2(load_address[5]), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_49), .A2(n_0_0_48), .ZN(n_0_0_41));
   NOR2_X1 i_0_0_142 (.A1(load_address[3]), .A2(load_address[2]), .ZN(n_0_0_42));
   OR4_X1 i_0_0_143 (.A1(load_address[12]), .A2(load_address[11]), .A3(
      load_address[10]), .A4(load_address[9]), .ZN(n_0_0_43));
   OR4_X1 i_0_0_144 (.A1(n_0_0_51), .A2(load_address[15]), .A3(load_address[14]), 
      .A4(load_address[13]), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_145 (.A1(load_address[1]), .A2(load_address[0]), .ZN(n_0_0_45));
   INV_X1 i_0_0_146 (.A(load_address[0]), .ZN(n_0_0_46));
   INV_X1 i_0_0_147 (.A(load_address[1]), .ZN(n_0_0_47));
   INV_X1 i_0_0_148 (.A(load_address[2]), .ZN(n_0_0_48));
   INV_X1 i_0_0_149 (.A(load_address[3]), .ZN(n_0_0_49));
   INV_X1 i_0_0_150 (.A(load_address[4]), .ZN(n_0_0_50));
   INV_X1 i_0_0_151 (.A(load_en), .ZN(n_0_0_51));
   INV_X1 i_0_0_152 (.A(reset), .ZN(n_0_0_52));
endmodule
